/* =====================================================================
    ____         _                 ____                      
   | __ )  _ __ (_)  __ _  _ __   / ___|  _   _  _ __    ___ 
   |  _ \ | '__|| | / _` || '_ \  \___ \ | | | || '_ \  / _ \
   | |_) || |   | || (_| || | | |  ___) || |_| || | | ||  __/
   |____/ |_|   |_| \__,_||_| |_| |____/  \__,_||_| |_| \___|
   
   =====================================================================
   Date: 2024-03
   Author: Brian Sune
   Contact: briansune@gmail.com
   Revision: 1.0.0
   FPGA: XC7A100FTG
   =====================================================================
*/

`timescale 1ns/1ps

module epp_basic(
	
	input wire					sys_clk_p,
	input wire					sys_clk_n,
	input wire					sys_nrst,
	
	input wire					btn_black,
	
	// clock gate driver
	output wire					epp_ckv,
	// gate start pulse
	output wire					epp_stv,
	// source output enable
	output wire					epp_xoe,
	// source start pulse
	output wire					epp_xstl,
	// source latch enable
	output wire					epp_xle,
	
	// clock source driver
	// SDCK = XCL - 33MHz
	output wire					epp_xcl,
	
	output wire					epp_mode,
	output wire		[7:0]		epp_data
);
	
	wire		epp_xcl_w;
	
	wire		glb_clk;
	wire		glb_nrst;
	
	clk_wiz_0 clk_inst0(
		.clk_out1	(glb_clk),
		.clk_out2	(epp_xcl_w),
		.locked		(glb_nrst),
		
		.resetn		(sys_nrst),
		.clk_in1_p	(sys_clk_p),
		.clk_in1_n	(sys_clk_n)
	);
	
	// in ns
	// localparam real ck_ns = 1000000000 / 20000000;
	// these parameters are minimum
	// localparam tle_dly		= 40;
	// localparam tle_w		= 150;
	// localparam tle_off		= 200;
	// =================================
	// make sure it is at least 1
	// localparam integer tle_dly_cyc	= (tle_dly / ck_ns) + 1;
	// localparam integer tle_w_cyc	= (tle_w / ck_ns) + 1;
	// localparam integer tle_off_cyc	= (tle_off / ck_ns) + 1;
	
	localparam lsl = 10;
	localparam lbl = 7;
	// 960 / [8 / 2bits]
	localparam ldl = 240;
	localparam lel = 105;
	localparam gdck_sta = 2;
	localparam gdck_hi = ldl * 2;
	localparam ltot = lsl + lbl + ldl + lel;
	
	localparam fsl = 1;
	localparam fbl = 4;
	localparam fdl = 540;
	localparam fel = 15;
	localparam ftot = fsl + fbl + fdl + fel;
	
	reg		[8 : 0]		cnt_a;
	reg		[10 : 0]	cnt_b;
	
	reg		[7 : 0]		epp_data_r;
	
	reg					sdle_r;
	reg					sdce_l_r;
	reg					gdck_r;
	
	reg					line_en;
	
	reg					gdsp_r;
	reg					sdoe_r;
	reg					gdoe_r;
	
	// reg					btn_black_r;
	
	assign epp_xcl		= epp_xcl_w;
	
	assign epp_xle		= sdle_r;
	
	assign epp_xoe		= sdoe_r;
	assign epp_mode		= gdoe_r;
	
	assign epp_ckv		= gdck_r;
	assign epp_xstl		= sdce_l_r;
	
	assign epp_stv		= gdsp_r;
	assign epp_data		= epp_data_r;
	
	reg		[2 : 0]		fsm_state;
	reg					run_load;
	reg					disp_all_w;
	reg					disp_all_b;
	reg		[3 : 0]		loop_cnt;
	
	reg		[4 : 0]		gray_cmp;
	
	localparam integer lut_bw = 20;
	
	reg		[lut_bw*2-1 : 0]	gray_lut	[0 : 15];
	
	initial begin
		// gray_lut[ 0] <= 24'b01_01_01_01_01_01_01_10_10_01_01_01;
		// gray_lut[ 1] <= 24'b00_01_01_01_01_01_01_01_10_10_01_01;
		// gray_lut[ 2] <= 24'b00_00_00_00_00_00_00_00_00_01_01_01;
		// gray_lut[ 3] <= 24'b00_00_00_00_00_00_00_00_00_00_01_01;
		// gray_lut[ 4] <= 24'b00_00_00_00_00_00_00_00_00_00_00_01;
		// gray_lut[ 5] <= 24'b00_00_00_10_10_10_10_10_01_01_01_01;
		// gray_lut[ 6] <= 24'b00_00_00_00_10_10_10_10_10_01_01_01;
		// gray_lut[ 7] <= 24'b00_00_00_00_00_10_10_10_10_10_01_01;
		// gray_lut[ 8] <= 24'b00_00_00_00_00_00_10_10_10_10_10_01;
		// gray_lut[ 9] <= 24'b00_00_00_00_01_01_01_01_01_01_01_10;
		// gray_lut[10] <= 24'b00_00_00_00_00_00_00_00_00_01_01_10;
		// gray_lut[11] <= 24'b00_00_00_00_01_01_01_01_01_01_10_10;
		// gray_lut[12] <= 24'b00_00_01_01_01_01_01_01_01_10_10_10;
		// gray_lut[13] <= 24'b00_01_01_01_01_01_01_01_10_10_10_10;
		// gray_lut[14] <= 24'b01_01_01_01_01_01_01_10_10_10_10_10;
		// gray_lut[15] <= 24'b00_00_00_00_00_00_00_10_10_10_10_10;
		
		gray_lut[ 0] <= 40'b01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01;
		gray_lut[ 1] <= 40'b01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_00;
		gray_lut[ 2] <= 40'b01_01_01_01_01_01_01_01_01_01_01_01_01_01_10_01_01_01_01_00;
		gray_lut[ 3] <= 40'b01_01_01_01_01_01_01_01_01_01_01_01_01_10_01_01_00_00_00_00;
		gray_lut[ 4] <= 40'b01_01_01_01_01_01_01_01_01_01_01_01_01_10_00_00_00_00_00_00;
		gray_lut[ 5] <= 40'b01_01_01_01_01_01_01_01_01_01_01_10_00_00_00_00_00_00_00_00;
		gray_lut[ 6] <= 40'b01_01_01_01_01_01_01_01_01_10_00_00_00_00_00_00_00_00_00_00;
		gray_lut[ 7] <= 40'b01_01_01_01_01_01_01_01_10_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[ 8] <= 40'b01_01_01_01_01_01_01_10_00_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[ 9] <= 40'b01_01_01_01_01_01_10_00_00_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[10] <= 40'b01_01_01_01_01_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[11] <= 40'b01_01_01_01_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[12] <= 40'b01_01_01_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[13] <= 40'b01_01_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[14] <= 40'b01_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;
		gray_lut[15] <= 40'b10_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;
	end
	
	// --------------------------------------
	localparam integer	fsm_reset		= 0,
						fsm_clean		= fsm_reset + 1,
						fsm_clean_loop	= fsm_clean + 1,
						fsm_draw		= fsm_clean_loop + 1,
						fsm_draw_wait	= fsm_draw + 1,
						fsm_done		= fsm_draw_wait + 1;
	// --------------------------------------
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			fsm_state <= fsm_reset;
			run_load <= 1'b0;
			disp_all_w <= 1'b0;
			disp_all_b <= 1'b0;
			loop_cnt <= 4'd0;
			gray_cmp <= 0;
		end else begin
			
			case(fsm_state)
				
				fsm_reset: begin
					run_load <= 1'b0;
					disp_all_w <= 1'b0;
					disp_all_b <= 1'b0;
					loop_cnt <= 4'd0;
					gray_cmp <= 0;
					
					fsm_state <= fsm_clean;
				end
					
				fsm_clean: begin
					if(loop_cnt < 4'd8)begin
						disp_all_b <= 1'b1;
						disp_all_w <= 1'b0;
					end else begin
						disp_all_b <= 1'b0;
						disp_all_w <= 1'b1;
					end
					
					run_load <= 1'b1;
					fsm_state <= fsm_clean_loop;
				end
				
				fsm_clean_loop: begin
					if(cnt_b >= (ftot - 1) && cnt_a >= (ltot - 1))begin
						run_load <= 1'b0;
						
						if(loop_cnt >= 4'd15)begin
							fsm_state <= fsm_draw;
							gray_cmp <= 0;
							loop_cnt <= 4'd0;
							disp_all_w <= 1'b0;
							disp_all_b <= 1'b0;
						end else begin
							fsm_state <= fsm_clean;
							loop_cnt <= loop_cnt + 1'b1;
						end
					end
				end
				
				fsm_draw: begin
					run_load <= 1'b1;
					fsm_state <= fsm_draw_wait;
				end
				
				fsm_draw_wait: begin
					if(cnt_b >= (ftot - 1) && cnt_a >= (ltot - 1))begin
						run_load <= 1'b0;
						
						if(gray_cmp >= (lut_bw-1) )begin
							fsm_state <= fsm_done;
							gray_cmp <= 0;
						end else begin
							fsm_state <= fsm_draw;
							gray_cmp <= gray_cmp + 1'b1;
						end
					end
				end
				
				fsm_done: begin
				
				end
				
				default: begin
					fsm_state <= fsm_clean;
					run_load <= 1'b0;
					disp_all_w <= 1'b0;
					disp_all_b <= 1'b0;
					loop_cnt <= 4'd0;
					gray_cmp <= 0;
				end
				
			endcase
		end
	end
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			cnt_a <= 9'd0;
		end else if(run_load)begin
			
			if(cnt_a >= (ltot - 1) )begin
				cnt_a <= 9'd0;
			end else begin
				cnt_a <= cnt_a + 1'b1;
			end
		end else begin
			cnt_a <= 9'd0;
		end
	end
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			cnt_b <= 11'd0;
		end else if(run_load)begin
			if(cnt_a >= (ltot - 1) )begin
				if(cnt_b >= (ftot - 1) )begin
					// cnt_b <= 11'd0;
				end else begin
					cnt_b <= cnt_b + 1'b1;
				end
			end
		end else begin
			cnt_b <= 11'd0;
		end
	end
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			sdle_r <= 1'b0;
		end else if(
			(cnt_b >= (fsl + fbl)) &&
			(cnt_b < (fsl + fbl + fdl))
		)begin
			if(cnt_a <= (lsl - 1) )begin
				sdle_r <= 1'b1;
			end else begin
				sdle_r <= 1'b0;
			end
		end else begin
			sdle_r <= 1'b0;
		end
	end
	
	// #####################################################
	// XSTL driver
	// #####################################################
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			sdce_l_r <= 1'b1;
		end else if(
			(cnt_b >= (fsl + fbl - 1)) &&
			(cnt_b < (fsl + fbl + fdl - 1))
		)begin
			if(
				(cnt_a >= (lsl + lbl - 1)) && 
				(cnt_a < (lsl + lbl + ldl - 1))
			)begin
				sdce_l_r <= 1'b0;
			end else begin
				sdce_l_r <= 1'b1;
			end
		end else begin
			sdce_l_r <= 1'b1;
		end
	end
	
	reg		[3839 : 0]		rom_data		[0 : 539];
	
	initial begin
		rom_data[0] <= 3840'h55555444444434333333333333233232323232323232323233223232232323232322322222223222222222222222222202000000000000000000000000000002022222234566555555556777655557CA7454445554324555555555444444444343333333332332323232323232232223222222223222222222322222222222222222222222222222222222222222222222222222222222222222222232222232222222222222222222222249CBBACCECCAABBBBCBBCCCCCCCCECCECECCCECCECECCBA7668ACCCCCCCCCAAEEECECECECECECBBBBBBCCA8554332355444444333332225432222222223222232322225555555555555444444434333333333333233232323232323232323233223232232323232322322222223222222222222222222202000000000000000000000000000002022222234566555555556777655557CA7454445554324555555555444444444343333333332332323232323232232223222222223222222222322222222222222222222222222222222222222222222222222222222222222222222232222232222222222222222222222249CBBACCECCAABBBBCBBCCCCCCCCECCECECCCECCECECCBA7668ACCCCCCCCCAAEEECECECECECECBBBBBBCCA855433235544444433333222543222222222322223232222;
		rom_data[1] <= 3840'h55544544444343333333333232332323232323232323232322333343332323223222223232322232323232323223232222000000000000000000000000000000022222335655555555555555555447BA63444455543345655545444544444343433333333233232322322322322223223223232322323232322232232323223222323232232222222222222222222232232232232323223232323232232223223232323232222222222202259AABCCCCCCBCCBCCCCCCCCCCCECCECCECEECEECCCECCC98788ABCCCCCCCACEECECCECECEEECCABBBCCCB8654333455544343333333235532223222322232222222225555555555544544444343333333333232332323232323232323232322333343332323223222223232322232323232323223232222000000000000000000000000000000022222335655555555555555555447BA63444455543345655545444544444343433333333233232322322322322223223223232322323232322232232323223222323232232222222222222222222232232232232323223232323232232223223232323232222222222202259AABCCCCCCBCCBCCCCCCCCCCCECCECCECEECEECCCECCC98788ABCCCCCCCACEECECCECECEEECCABBBCCCB865433345554434333333323553222322232223222222222;
		rom_data[2] <= 3840'h555545444444333433333333333232322322322323232322345555555343443323232323222232222223222223222222322000000200000000000000000000000002234455555554554444454544479854443455554236776555545444434434343333233323232232232232232322322322222232222222223222222222222222222222222222232223222322232222222222222222222222222223232322322222222222322222222222238BBBBCCCCCCCCCCCCCCCCBBCCCCCCECEECEECCEECECECB98878ACCECECCCEEECECECECECEEEBABCECEC975553325554334333333333365322222322232223232232255555555555545444444333433333333333232322322322323232322345555555343443323232323222232222223222223222222322000000200000000000000000000000002234455555554554444454544479854443455554236776555545444434434343333233323232232232232232322322322222232222222223222222222222222222222222222232223222322232222222222222222222222222223232322322222222222322222222222238BBBBCCCCCCCCCCCCCCCCBBCCCCCCECEECEECCEECECECB98878ACCECECCCEEECECECECECEEEBABCECEC9755533255543343333333333653222223222322232322322;
		rom_data[3] <= 3840'h555554444443434333333323223232223233333232334444567777665555554432222223223222322322232222232232322200000220000000000000000000000020233333444444443344444444457644443334553235778865444444444343343333333332322222322322322322223222322222232232232223222322232222232222322232222222222222222222222222222232223223223222222222222322322322222222222222225ACABCCEECCCCCCCECCCCCCCCCCCCECEEEECEECCCECCCCA87778BCECCCEEEECCECECECEECEBBBBCCEEC876553335543332223333333367532222223222222222222255555555555554444443434333333323223232223233333232334444567777665555554432222223223222322322232222232232322200000220000000000000000000000020233333444444443344444444457644443334553235778865444444444343343333333332322222322322322322223222322222232232232223222322232222232222322232222222222222222222222222222232223223223222222222222322322322222222222222225ACABCCEECCCCCCCECCCCCCCCCCCCECEEEECEECCCECCCCA87778BCECCCEEEECCECECECEECEBBBBCCEEC8765533355433322233333333675322222232222222222222;
		rom_data[4] <= 3840'h5555545444443333333333323323233323345554344556678888777765567755443333222222222222222222222222222222000000000000000000000000000000002223233333333433334343443454445333355432245789865444444344343333333323232322322322322222223222222232222222222222222222222222322222222222222222222322232222322232222322222222222222232322222222222222232232222222222236AACCCCCECECCCCCCCCCCCCCECEECEECECECCCCCCCCCBA976789BCEEEEEECECCECECECECCBBCCCCECA8765543453322222222233333687533222222222322222222555555555555545444443333333333323323233323345554344556678888777765567755443333222222222222222222222222222222000000000000000000000000000000002223233333333433334343443454445333355432245789865444444344343333333323232322322322322222223222222232222222222222222222222222322222222222222222222322232222322232222322222222222222232322222222222222232232222222222236AACCCCCECECCCCCCCCCCCCCECEECEECECECCCCCCCCCBA976789BCEEEEEECECCECECECECCBBCCCCECA8765543453322222222233333687533222222222322222222;
		rom_data[5] <= 3840'h555545444443433433333334334334444456777665678888999876666566655554444332232232232232322232222222232202000000000000000000000000000000020222222223333343333333322334343335543233567887654444444343333333333232322322322222232232222232222222222322222322222222222222232222222222222222222222222222222222222222222222222222222232222222222222222232222222222358ABCCCCCCCEECECECCCCECCEECEECECCCECCCCCCCCAA987789CCEEEEEEECECECECECCCCBBCCBBBA9876553355422222222222233378776522222232222222222255555555555545444443433433333334334334444456777665678888999876666566655554444332232232232232322232222222232202000000000000000000000000000000020222222223333343333333322334343335543233567887654444444343333333333232322322322222232232222232222222222322222322222222222222232222222222222222222222222222222222222222222222222222222232222222222222222232222222222358ABCCCCCCCEECECECCCCECCEECEECECCCECCCCCCCCAA987789CCEEEEEEECECECECECCCCBBCCBBBA98765533554222222222222333787765222222322222222222;
		rom_data[6] <= 3840'h55554555444334333333345555555555555777888888889999876777656765545555555433333322322222322232223222222020000000000000000000000000000000202222222222233332333233223333334454443346667776544343434333333332332322322222222322222222222222232232222232222223222222222222222222222222222222222222322232222222222222222223223223222222232223223223222222222222222478ABCCCCCCCCCCCECEECEECEECEECCECCCCCCCCCCAAA98889BCCEEEECCCCCCCECECECCBCBBBAAA887755446533323333322022336755663222222222222222225555555555554555444334333333345555555555555777888888889999876777656765545555555433333322322222322232223222222020000000000000000000000000000000202222222222233332333233223333334454443346667776544343434333333332332322322222222322222222222222232232222232222223222222222222222222222222222222222222322232222222222222222223223223222222232223223223222222222222222478ABCCCCCCCCCCCECEECEECEECEECCECCCCCCCCCCAAA98889BCCEEEECCCCCCCECECECCBCBBBAAA88775544653332333332202233675566322222222222222222;
		rom_data[7] <= 3840'h55555544444434344544456766667777776777888988888998877787777776544445555554544433222222222222222222222222020000000000000000000000000000202022022222222222222333233432333434555545556777755443433333333233323223223223223223222322322232222222232222222222222222222222222222222222222222222222222222232222222222222222222222222232222222222222222222222222222258ABBCCCECCCCCECCECEEEECECECECECEECECECCCCCCBB989ABCEEEEECECECECECECCCCCCBBAA9988755556432222333333223225654443222222222222222225555555555555544444434344544456766667777776777888988888998877787777776544445555554544433222222222222222222222222020000000000000000000000000000202022022222222222222333233432333434555545556777755443433333333233323223223223223223222322322232222222232222222222222222222222222222222222222222222222222222232222222222222222222222222232222222222222222222222222222258ABBCCCECCCCCECCECEEEECECECECECEECECECCCCCCBB989ABCEEEEECECECECECECCCCCCBBAA998875555643222233333322322565444322222222222222222;
		rom_data[8] <= 3840'h5555454444445556676566777677778777767788899888899987888877888775433344445445555443223222222222222222222222220000000000000000000000000220220220222222222222233322475434432345554455577787754333433333332323232222232222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222223222222222322322222232222232222223589ABECCCCCBBBECCECEEEEEECECECCCECCEEECCECCCB9888ACEEEEEECCCECECEEECCCBAABBBA98876555532200222222222322455533222222222222222222555555555555454444445556676566777677778777767788899888899987888877888775433344445445555443223222222222222222222222220000000000000000000000000220220220222222222222233322475434432345554455577787754333433333332323232222232222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222223222222222322322222232222232222223589ABECCCCCBBBECCECEEEEEECECECCCECCEEECCECCCB9888ACEEEEEECCCECECEEECCCBAABBBA98876555532200222222222322455533222222222222222222;
		rom_data[9] <= 3840'h55555445556667888887767766678887777778888988889A99888888788887765333333333334555543222222222232222222222222222000000000000000000000002022022020220222020222222323653467432233544556788899864433333333232323223222222222222222222222222322222222222222222222222222222222222222222222222222222223222222222222222222222222222222222222322222223222222222222222222457ABBCBB99ABCCCCEECEEEEEECCCCCCCCECCCCCCCBBA8889ACEEEEECECCECEECECCBA9ABCBA988766655422222202020022224654332222222222222222225655555555555445556667888887767766678887777778888988889A99888888788887765333333333334555543222222222232222222222222222000000000000000000000002022022020220222020222222323653467432233544556788899864433333333232323223222222222222222222222222322222222222222222222222222222222222222222222222222222223222222222222222222222222222222222222322222223222222222222222222457ABBCBB99ABCCCCEECEEEEEECCCCCCCCECCCCCCCBBA8889ACEEEEECECCECEECECCBA9ABCBA98876665542222220202002222465433222222222222222222;
		rom_data[10] <= 3840'h55555556789999989988767766788889888889AAA99899AAA9888888788888776543222322333345554443333332222222222222222222222000000000000000000000220000202020202022020222222322355422223454555689AABA976543323233323223222222223222322222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222223222223222222222222259AABBA99ACCCCEEEEEEECCEECECECECCCCCCCCBBBA998AABEEEEEECCCCCCEECCCBAABCCBAA98776545443333322222202235754333222222222222222226555555555555556789999989988767766788889888889AAA99899AAA9888888788888776543222322333345554443333332222222222222222222222000000000000000000000220000202020202022020222222322355422223454555689AABA976543323233323223222222223222322222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222223222223222222222222259AABBA99ACCCCEEEEEEECCEECECECECCCCCCCCBBBA998AABEEEEEECCCCCCEECCCBAABCCBAA9877654544333332222220223575433322222222222222222;
		rom_data[11] <= 3840'h555667789BCCCBA9988776778888999999999BBBBA999BBA987788877888888875533232232323345555554445432222222222222222222220200000000000000000000000000020020202202020220000022322223344455556799AABA988755332323232222232222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222232222223222222222222222479AA9AAABCBCEEEEEECEEEECECCECECCECCCCCCBBBAAA999CEEEEEECECECECCCCBBBCCCBBA988775554444333333322233346533332222222222222222256555555555667789BCCCBA9988776778888999999999BBBBA999BBA987788877888888875533232232323345555554445432222222222222222222220200000000000000000000000000020020202202020220000022322223344455556799AABA988755332323232222232222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222232222223222222222222222479AA9AAABCBCEEEEEECEEEECECCECECCECCCCCCBBBAAA999CEEEEEECECECECCCCBBBCCCBBA9887755544443333333222333465333322222222222222222;
		rom_data[12] <= 3840'h5568888ACCEECCB9888776789999999AA99AAABBBAAAABBA97777776778887788754333232232333345555555555433222222222222222222222200000000000000000000000000200202002000002000020222022344444455567899998888875333223232322232222222222222222222222222222222222222222222222222222222222222222222222222222222322222222222222222222222222222222222232222222222222222222222222222356579AAAABCCCCECEECEEEEEEECECCECCECCCCBBCBBA989AEEEEEECCCCECCCBBBBCECCBBA9988755543443334333453343355324432222222222222222655555555568888ACCEECCB9888776789999999AA99AAABBBAAAABBA97777776778887788754333232232333345555555555433222222222222222222222200000000000000000000000000200202002000002000020222022344444455567899998888875333223232322232222222222222222222222222222222222222222222222222222222222222222222222222222222322222222222222222222222222222222222232222222222222222222222222222356579AAAABCCCCECEECEEEEEEECECCECCECCCCBBCBBA989AEEEEEECCCCECCCBBBBCECCBBA9988755543443334333453343355324432222222222222222;
		rom_data[13] <= 3840'h677899ACEEEEEEC9888777899A9999A999A9ABAAAAAAABBA876566555676666777755433322232233334444555555432222222222222222222222222000000000000000000000000002000200002000000002020223333334455558888877789985533322222222222222222222222222222222222222222222222222222222222222222222022222222222222222222222222222222222222222222222222222222222222232222223222222222222222222457899BCCCCECECEECECCEECECECECCCCBBBEECCB999AACEEEEEECECECBAABCCCCCCBAA98875544333343333455434335520232222222222222222255555556677899ACEEEEEEC9888777899A9999A999A9ABAAAAAAABBA876566555676666777755433322232233334444555555432222222222222222222222222000000000000000000000000002000200002000000002020223333334455558888877789985533322222222222222222222222222222222222222222222222222222222222222222222022222222222222222222222222222222222222222222222222222222222222232222223222222222222222222457899BCCCCECECEECECCEECECECECCCCBBBEECCB999AACEEEEEECECECBAABCCCCCCBAA988755443333433334554343355202322222222222222222;
		rom_data[14] <= 3840'h8889ABCCEEEEEECB98877899AAAA9A9AA9A9AA9999999AAA887655555555555777775554332232323333333334445543322222222222222222222222220000000000000000000000000020000020000000000020223333233333456777777778999885432222222222222222222222222222222222222222222222022022022222222222222222222222222222222222222222222222222222222222222222222222222232222232222222222222222222222223578ABBCCCCCCCCECECCECECECCECCBBCEEEECCBA99BCEEEEEECECCCBAABCEECCCBAA998644433433334333444454355220222222222222222222666677878889ABCCEEEEEECB98877899AAAA9A9AA9A9AA9999999AAA887655555555555777775554332232323333333334445543322222222222222222222222220000000000000000000000000020000020000000000020223333233333456777777778999885432222222222222222222222222222222222222222222222022022022222222222222222222222222222222222222222222222222222222222222222222222222232222232222222222222222222222223578ABBCCCCCCCCECECCECECECCECCBBCEEEECCBA99BCEEEEEECECCCBAABCEECCCBAA998644433433334333444454355220222222222222222222;
		rom_data[15] <= 3840'h99ABBBCEEEEEECCBA88889ABBAAA9AA9999A98888899998988765555666554567777666554333333333333333334444433222222222222222222222222222000000000000000000000000000022200000000000022333322223445557666777889ABB98542222222222222222222222222222222222222222222222222222220220202022022222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222479AAABBBBCEEEEECECEECCCEBBBCEEEECCCCCBB9ABCEEEEEEECEBBBBCCCCCCCBBA9975533344433333333344544443222222222222222222227789999A99ABBBCEEEEEECCBA88889ABBAAA9AA9999A98888899998988765555666554567777666554333333333333333334444433222222222222222222222222222000000000000000000000000000022200000000000022333322223445557666777889ABB98542222222222222222222222222222222222222222222222222222220220202022022222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222479AAABBBBCEEEEECECEECCCEBBBCEEEECCCCCBB9ABCEEEEEEECEBBBBCCCCCCCBBA997553334443333333334454444322222222222222222222;
		rom_data[16] <= 3840'hBBBCCEEEEEEEEECBB99899BBBAAAAAAA9999877778889888888755677777555577777666554334333323333334433344433333222222222220222022222222200000000000000000000000000020000000000000223333223334555555566778889ACCCC86432222222222222222222222222222222222222222222202222222222222222220222222222222222222222222222222222222222222222222222222222222222232222222222222222222222222022259B9989ABCCCECECCEEEEEECBCCCCCAAAAABECCBA9BEEEEEEEECBBBBCECEECCBBAA964454554444423333344444443222222222222222222229AAABBCBBBBCCEEEEEEEEECBB99899BBBAAAAAAA9999877778889888888755677777555577777666554334333323333334433344433333222222222220222022222222200000000000000000000000000020000000000000223333223334555555566778889ACCCC86432222222222222222222222222222222222222222222202222222222222222220222222222222222222222222222222222222222222222222222222222222222232222222222222222222222222022259B9989ABCCCECECCEEEEEECBCCCCCAAAAABECCBA9BEEEEEEEECBBBBCECEECCBBAA96445455444442333334444444322222222222222222222;
		rom_data[17] <= 3840'hCBCCEEEEEEEEECECBAA99ABBBAAA9A9999988666788889888887667788875556777777766555555433333333344443444444443222222220222222222222222220000000000000000000000000000000000000000223332333343445555557777789ABEEECA87532222222222222222222222222222220222222022222022022222222222222222222222222222222222223222222222222222222222222222222222223222222232222222222222222202202222236887788AB86566689ABCCCA9AAA999999AABCEC98ACEEEEEEECCCCCCECCCCCCBBB86445576444443444345555554222222222222222222222CCCCCCCCCBCCEEEEEEEEECECBAA99ABBBAAA9A9999988666788889888887667788875556777777766555555433333333344443444444443222222220222222222222222220000000000000000000000000000000000000000223332333343445555557777789ABEEECA87532222222222222222222222222222220222222022222022022222222222222222222222222222222222223222222222222222222222222222222222223222222232222222222222222202202222236887788AB86566689ABCCCA9AAA999999AABCEC98ACEEEEEEECCCCCCECCCCCCBBB86445576444443444345555554222222222222222222222;
		rom_data[18] <= 3840'hCCCCEEEEEECECECCBBAAAAAAAA9999999889865677788998888766778887555677788777655556543223233334343434344555532222022222222222022222222220000000000000000000000000000000000000222232223332334556555567778899ABECECCA87532222222222222222222222222222222022220222222222022022022022202222222222222222222222222222222222222222222222222222222222222222223222222222222222222222220223343357985222334556788778888889899ABCEEB99AACEEEEEECCCCECECECCCCBB95445555445434454333455554222222222222222222222EEEEEEECCCCCEEEEEECECECCBBAAAAAAAA9999999889865677788998888766778887555677788777655556543223233334343434344555532222022222222222022222222220000000000000000000000000000000000000222232223332334556555567778899ABECECCA87532222222222222222222222222222222022220222222222022022022022202222222222222222222222222222222222222222222222222222222222222222223222222222222222222222220223343357985222334556788778888889899ABCEEB99AACEEEEEECCCCECECECCCCBB95445555445434454333455554222222222222222222222;
		rom_data[19] <= 3840'hCCCEEEEECCCCCCCCCCBBAAA9A998899988988766777789998887777777755556778888876555675432323323433333344444444433222222222022222220222222220000000000000000000000000000000000002222222233323345555545577888889AABBCCCCB975320202020202020202220220222222222222202220222222222222222222222222222222222222222222222222222222222222222222222222322232223222222222222222222222222222222222224753222333455556677888ABBCCCEEEEEEBA9ACEEEEEEEA9A9CCECCECCBC84445554455444454333444454322222222222222222222EEEECECECCCEEEEECCCCCCCCCCBBAAA9A998899988988766777789998887777777755556778888876555675432323323433333344444444433222222222022222220222222220000000000000000000000000000000000002222222233323345555545577888889AABBCCCCB975320202020202020202220220222222222222202220222222222222222222222222222222222222222222222222222222222222222222222222322232223222222222222222222222222222222222224753222333455556677888ABBCCCEEEEEEBA9ACEEEEEEEA9A9CCECCECCBC84445554455444454333444454322222222222222222222;
		rom_data[20] <= 3840'hECCCCEECBBBBCCCCCCCBBAAA998888888899887777778888988776666665555667888877766566543333333333334334443333344322222220222202022220220222220000000000000000000000000020000000202020222323344445555556677778888889ABBCCA86543222202222222202222222220222220222220222202202202202222222222222222222222222222222222222222222222222222222222222222223222222232222222222222022022222022020223322223334454479CCCCEEEEEEEEEEEEEEBABBEEEEEEE97779BCEECCCCB74344433454334544445443443222222222222222222222EEEEEEECECCCCEECBBBBCCCCCCCBBAAA998888888899887777778888988776666665555667888877766566543333333333334334443333344322222220222202022220220222220000000000000000000000000020000000202020222323344445555556677778888889ABBCCA86543222202222222202222222220222220222220222202202202202222222222222222222222222222222222222222222222222222222222222222223222222232222222222222022022222022020223322223334454479CCCCEEEEEEEEEEEEEEBABBEEEEEEE97779BCEECCCCB74344433454334544445443443222222222222222222222;
		rom_data[21] <= 3840'hCCCCCECCBAABCCCCECCCBBBAA99888888899888888777888898876666555567667788887777766655433333444344344434333344443202222222222222222222222222000000000000000000000000002000002020000222222343334455555545577877668899ABCBBB887543222222222222222220222202222222222222222222222222022222222222222222222222222222222222222222222222222222222222222222223232222222222222222222202222202222022222233334558CEEEEEEEEEEEEEEEEEEEECB9AEEEEEEA87778BECECCEA53324323443344555444444444322222222222222222222EEECCCCCCCCCCECCBAABCCCCECCCBBBAA99888888899888888777888898876666555567667788887777766655433333444344344434333344443202222222222222222222222222000000000000000000000000002000002020000222222343334455555545577877668899ABCBBB887543222222222222222220222202222222222222222222222222022222222222222222222222222222222222222222222222222222222222222222223232222222222222222222202222202222022222233334558CEEEEEEEEEEEEEEEEEEEECB9AEEEEEEA87778BECECCEA53324323443344555444444444322222222222222222222;
		rom_data[22] <= 3840'hBABBBCBBBABBBBCCCCCBBBBBBB99888888899888877778888888876665556777677889887877776655433333434334334333333445543220222020222022022220222222000000000000000000000000200000002000000022022333334455543345567755689AAAAABBBAABBA75532222022202202222222222022022020202202202202222222222222222222222222222222222222222222222222222222222222223222222222222222222222222220222222022222022020222223479CEEEEEEEEEEEEEEEEEEEEEEEB86CEEEEEB987779CECECE953323333433444344433435444422222222222222222222ECECECCBBABBBCBBBABBBBCCCCCBBBBBBB99888888899888877778888888876665556777677889887877776655433333434334334333333445543220222020222022022220222222000000000000000000000000200000002000000022022333334455543345567755689AAAAABBBAABBA75532222022202202222222222022022020202202202202222222222222222222222222222222222222222222222222222222222222223222222222222222222222222220222222022222022020222223479CEEEEEEEEEEEEEEEEEEEEEEEB86CEEEEEB987779CECECE953323333433444344433435444422222222222222222222;
		rom_data[23] <= 3840'hAAAAABAABBBBAABCCCBBBBBBBBAA88888889888887777788888887776556677667789898888887766654333433343333334333345555322220222220222222202222222222000000000000020000000020000000000000022020222333334443334455655579BBA87766667898998875422220222222220222222202222222222222222220222022222222222222222222222222222222222222222222222222222222222223222222222222222222220222222222202222202222222225BEEEEEEEEEEEEEEEEEEEEEEEEEE937CEEEEE987778ACEECC733333343444433333333334422332222222222222222222CECCCCCBAAAAABAABBBBAABCCCBBBBBBBBAA88888889888887777788888887776556677667789898888887766654333433343333334333345555322220222220222222202222222222000000000000020000000020000000000000022020222333334443334455655579BBA87766667898998875422220222222220222222202222222222222222220222022222222222222222222222222222222222222222222222222222222222223222222222222222222220222222222202222202222222225BEEEEEEEEEEEEEEEEEEEEEEEEEE937CEEEEE987778ACEECC733333343444433333333334422332222222222222222222;
		rom_data[24] <= 3840'hA999AABBABBBAABBCBBBBBBBBBBA99889888888777777888888778777555666667888988888888776654323333334333343334445675432222022022222220222222222222222000000000000000000000000000000000002222222233334433334555556678985432223334444689A9875432220222022220202222220220220220220222222222222222222222222322222222222222222222222222222222222223222222232232222222222222222222202202222020220202222349EEEEEEEEEEEEEEEEEEEEEEEEEEEB23AEEEEEC8667678BCEB532333443454433333333223322232222222222222222222CCCECCBBA999AABBABBBAABBCBBBBBBBBBBA99889888888777777888888778777555666667888988888888776654323333334333343334445675432222022022222220222222222222222000000000000000000000000000000000002222222233334433334555556678985432223334444689A9875432220222022220202222220220220220220222222222222222222222222322222222222222222222222222222222222223222222232232222222222222222222202202222020220202222349EEEEEEEEEEEEEEEEEEEEEEEEEEEB23AEEEEEC8667678BCEB532333443454433333333223322232222222222222222222;
		rom_data[25] <= 3840'hBAAAAAAABBBBAAABBBBBBBAAAAAA99998888887777888888888777777555656777889999888888877654332333344333544345556786543222220222020202222022022222220000000000000000000000000000000000000202222233333333344455556675532220002202233246899AA9764322202222222222202222222022022022222222222222222222222322222222222222222222222222222222222222222232222222222222222222222220220220222222220202220259EEEEEEECCEECC99ACEEEEEEEEEEEEC227EEEEEE865554579C8422323343443333443333333320222222222222222222222CCCCCCCBBAAAAAAABBBBAAABBBBBBBAAAAAA99998888887777888888888777777555656777889999888888877654332333344333544345556786543222220222020202222022022222220000000000000000000000000000000000000202222233333333344455556675532220002202233246899AA9764322202222222222202222222022022022222222222222222222222322222222222222222222222222222222222222222232222222222222222222222220220220222222220202220259EEEEEEECCEECC99ACEEEEEEEEEEEEC227EEEEEE865554579C8422323343443333443333333320222222222222222222222;
		rom_data[26] <= 3840'hBBBBAAABABAAAAAAABAAAAAAAAA999899888788878878888888776777765556677889999898888887765433223455335665457788887553302022202222222202222222222222000000000000000000000000000000000000000222222333323333445555543232202000000022222479BCCA875543222020222022220220222222222222022022222222222222222222222222222222222222222222222222222222222223222222222222222222222222222222220220220220225CEEEEEEC99A9988778AABECECCECEEEC4039EEEEEABA75557885232334323343334344443333320222222222222222222222CCCCCCCBBBBBAAABABAAAAAAABAAAAAAAAA999899888788878878888888776777765556677889999898888887765433223455335665457788887553302022202222222202222222222222000000000000000000000000000000000000000222222333323333445555543232202000000022222479BCCA875543222020222022220220222222222222022022222222222222222222222222222222222222222222222222222222222223222222222222222222222222222222220220220220225CEEEEEEC99A9988778AABECECCECEEEC4039EEEEEABA75557885232334323343334344443333320222222222222222222222;
		rom_data[27] <= 3840'hBCBBBBBABBABBA9AAAA9AA9AAA9999988888878788787888888877778776566678899999998889888766543322455345677788888987555432220222020220222202222222222000000000000000000000000000000000000000020222222223233344454322234202233322222202235688777778864322220222222222220202202020222222222222222222222223222222222222222222222022222222222222232222222222322222222222222202222020220222220220228CEEEEEEC988877666787888ABCCBBBBCC83248EEE958865677753223333333334344333333333322222222222222222222222CCCCBCBBBCBBBBBABBABBA9AAAA9AA9AAA9999988888878788787888888877778776566678899999998889888766543322455345677788888987555432220222020220222202222222222000000000000000000000000000000000000000020222222223233344454322234202233322222202235688777778864322220222222222220202202020222222222222222222222223222222222222222222222022222222222222232222222222322222222222222202222020220222220220228CEEEEEEC988877666787888ABCCBBBBCC83248EEE958865677753223333333334344333333333322222222222222222222222;
		rom_data[28] <= 3840'hCCCBBBBABABBAAAAAAA999A9A9A999998887888787877788887877778876665678888999998889988776553323344445678899988885545554322202222022222222202222220000000000000000000000000000000000000000002002020222323333343200244433455553345532222223224789AA875422202022022022222022222222222222222222222222222222222222222222222222222222222222222222223222232222223222222222222222222202222202222024CEEEEECA9987877778887566788889AA9AB8522698644455555433223323343333333334333333443222222222222222222222CCBCCCBCCCCBBBBABABBAAAAAAA999A9A9A999998887888787877788887877778876665678888999998889988776553323344445678899988885545554322202222022222222202222220000000000000000000000000000000000000000002002020222323333343200244433455553345532222223224789AA875422202022022022222022222222222222222222222222222222222222222222222222222222222222222222223222232222223222222222222222222202222202222024CEEEEECA9987877778887566788889AA9AB8522698644455555433223323343333333334333333443222222222222222222222;
		rom_data[29] <= 3840'hCCCCBBBABBBBBAAAAAA9999A9A9A9998877777778777778888777778887765568888899AA9888998888765433233444557889A9888654455555320220222202020220222222000000000000000000000000000000000000000000000200202022222223320022334444445555576655430000004788A9AA975332202222220222222020202202222222222222222222222222222222222222222222222222222222222222223222222322222222222222202222222020222020249EEEEEB9888778888999877667777778889ACB74245553334444322233233333332222235554434544322222222222222222222CCCCCBCBCCCCBBBABBBBBAAAAAA9999A9A9A9998877777778777778888777778887765568888899AA9888998888765433233444557889A9888654455555320220222202020220222222000000000000000000000000000000000000000000000200202022222223320022334444445555576655430000004788A9AA975332202222220222222020202202222222222222222222222222222222222222222222222222222222222222223222222322222222222222202222222020222020249EEEEEB9888778888999877667777778889ACB74245553334444322233233333332222235554434544322222222222222222222;
		rom_data[30] <= 3840'hBCCCCBBAAABBBBBBBAA999999A9AA99888778887777777788877788888775557888888AAA9999999888877543333355557889A9987554444555542022020222222222222220000000000000000000000000000000000000000000000000002022222233322022233333345555555555543000002578888ACCA8754320000220202022222222222222222222222222222222222222222222222222222222222222222222322222223222222222222222222222202222220222023AEEEEEA8877778899899999999988877799ACCEC8222333333332222333322335557885434567754444322222222222222222222CCCCCCBBBCCCCBBAAABBBBBBBAA999999A9AA99888778887777777788877788888775557888888AAA9999999888877543333355557889A9987554444555542022020222222222222220000000000000000000000000000000000000000000000000002022222233322022233333345555555555543000002578888ACCA8754320000220202022222222222222222222222222222222222222222222222222222222222222222222322222223222222222222222222222202222220222023AEEEEEA8877778899899999999988877799ACCEC8222333333332222333322335557885434567754444322222222222222222222;
		rom_data[31] <= 3840'hCBBCBBBA9ABBBCBBBBA988899A9AA989888888877777777888888999888755578898889A9999AAA98999887544334687778889988775445445555322022220202202222220200000000000000000000000000000000000000000000000000000002023332222223323334555443333344432322246876789BCCCBA754432202222222022022222222222222222222222222222222222222222222222222222222222222222222222222232222222222202220222022222222227EEEEEB987776788888888AAAAB9A9A988ACCCCBB8400002222222002333222336769EEC876446765333332222222222222222222CCCCCBBBCBBCBBBA9ABBBCBBBBA988899A9AA989888888877777777888888999888755578898889A9999AAA98999887544334687778889988775445445555322022220202202222220200000000000000000000000000000000000000000000000000000002023332222223323334555443333344432322246876789BCCCBA754432202222222022022222222222222222222222222222222222222222222222222222222222222222222222222232222222222202220222022222222227EEEEEB987776788888888AAAAB9A9A988ACCCCBB8400002222222002333222336769EEC876446765333332222222222222222222;
		rom_data[32] <= 3840'hBBBBBBAAAAACBCCCBBB9988999AA99898887888777777777888899A9888765568888899999899A9999A9887655545787777889A9987544555455553220202222022220202220000000000000000000000000000000000000000000000000000000022332022223233333344443332333332222235677677889ABCCECEB8754222020220222222202222222222222222222222222222222222222222222222222222222232232232223222232222222222222222220202222025BEEEAA98877778888877878888989A98877ACA9995300000000000022233233455546989CEC842355422222222222222222222222CBBCBBBCBBBBBBAAAAACBCCCBBB9988999AA99898887888777777777888899A9888765568888899999899A9999A9887655545787777889A9987544555455553220202222022220202220000000000000000000000000000000000000000000000000000000022332022223233333344443332333332222235677677889ABCCECEB8754222020220222222202222222222222222222222222222222222222222222222222222222232232232223222232222222222222222220202222025BEEEAA98877778888877878888989A98877ACA9995300000000000022233233455546989CEC842355422222222222222222222222;
		rom_data[33] <= 3840'hBBBBBBABAABBCCBCCBBA988999AAA9888878888777788877788999A998877657788889A988899A9A9AA988876654478878888AAAA9865455555565422202202022020222222220000000000000000000000000000000000000000000000000000020033200222222332222343222232332202223565567878889BCCEEEEEEA874322202202222222222222222222222222222222222222222222222222222222222322322222222222222222222222222220202222222022037BBA88888877788998777655556767767877999AB96320000000000022233347777778988BAAB85332333222222222222222222222CCCBBBBBBBBBBBABAABBCCBCCBBA988999AAA9888878888777788877788999A998877657788889A988899A9A9AA988876654478878888AAAA9865455555565422202202022020222222220000000000000000000000000000000000000000000000000000020033200222222332222343222232332202223565567878889BCCEEEEEEA874322202202222222222222222222222222222222222222222222222222222222222322322222222222222222222222222220202222222022037BBA88888877788998777655556767767877999AB96320000000000022233347777778988BAAB85332333222222222222222222222;
		rom_data[34] <= 3840'hBBBAAAAAAABBBBCBBBBA99899AABA9898888888878888877788899999887777778888999988999A99A98898876555788888899AAA98755555555665322020222222222222202222332000000000000000000000000000000000000000000000000020233002222222200022222202232220000235555777768889BCCEEEEEEEECA8432022202022222222222222222222222222222222222222220222222222222222222322322232222322222222222222222220220222237BB898888887689998875555555555457ACA99999864320000000000002236755555776778BA9AEC730243222222222222222222222CCBBBCBBBBBAAAAAAABBBBCBBBBA99899AABA9898888888878888877788899999887777778888999988999A99A98898876555788888899AAA98755555555665322020222222222222202222332000000000000000000000000000000000000000000000000020233002222222200022222202232220000235555777768889BCCEEEEEEEECA8432022202022222222222222222222222222222222222222220222222222222222222322322232222322222222222222222220220222237BB898888887689998875555555555457ACA99999864320000000000002236755555776778BA9AEC730243222222222222222222222;
		rom_data[35] <= 3840'hBBBAABAAAAAABBBBBBBA9889ABBAA998888888887888887788898999988877778887899888899A9AA999999987557888888898AA9888654555555654222222020202022022222224432000000000000000000000000000000000000000000000000003530202220000000002222222222202223334555676778889ACCCEEEEEEEEEE8532202222222222222222222222322222222222222222222222222222222222322222322222232222322222222202222022220222027CCB99888887779BA8876555555555447BEEB8555544430000000000002223543454567655579ABBCE82243222222222222222222222CCCCCBCBBBBAABAAAAAABBBBBBBA9889ABBAA998888888887888887788898999988877778887899888899A9AA999999987557888888898AA9888654555555654222222020202022022222224432000000000000000000000000000000000000000000000000003530202220000000002222222222202223334555676778889ACCCEEEEEEEEEE8532202222222222222222222222322222222222222222222222222222222222322222322222232222322222222202222022220222027CCB99888887779BA8876555555555447BEEB8555544430000000000002223543454567655579ABBCE82243222222222222222222222;
		rom_data[36] <= 3840'hCBBBBAAA9AAAABBBABA99999ABBA999888888888889888878888999A998777777778889888889A9AAAA999A987767888888999AA9888655555555564320202222222222222222223330000000000000000000000000000000000000000000000000002440000202000000220223542222232322234544567777788ACEECEEEEEEEEEEBA7543222020222222222222322222322232222222222222222222222222222222232222232222322223222222222022220222222249B9A99888777778B9887545555555445AEEC95323444542000000000002223345555689778ACAABCA993243222222222222222222222ECCCCCCCCBBBBAAA9AAAABBBABA99999ABBA999888888888889888878888999A998777777778889888889A9AAAA999A987767888888999AA9888655555555564320202222222222222222223330000000000000000000000000000000000000000000000000002440000202000000220223542222232322234544567777788ACEECEEEEEEEEEEBA7543222020222222222222322222322232222222222222222222222222222222232222232222322223222222222022220222222249B9A99888777778B9887545555555445AEEC95323444542000000000002223345555689778ACAABCA993243222222222222222222222;
		rom_data[37] <= 3840'hCCCCCBBAAAAAAA9AAA998899BAAA998888888888889888878899999A99877777777888888889999AAA9AAAA998877878888999A998987655655545553220220202020220220222223220000000000000000000000000000000000000000000000000022200002000000033222248522023333223344455576667778BCCECCEEEEEEEEECCB9875433322222222222222222222222223222222222222222222222222232222232322232222222222222222222222222020226BA899888877787789875455555554448EECC832224444330000000000002355556776788888ABBEEB874023222222222222222222222EEEECECCCCCCCBBAAAAAAA9AAA998899BAAA998888888888889888878899999A99877777777888888889999AAA9AAAA998877878888999A998987655655545553220220202020220220222223220000000000000000000000000000000000000000000000000022200002000000033222248522023333223344455576667778BCCECCEEEEEEEEECCB9875433322222222222222222222222223222222222222222222222222232222232322232222222222222222222222222020226BA899888877787789875455555554448EECC832224444330000000000002355556776788888ABBEEB874023222222222222222222222;
		rom_data[38] <= 3840'hCCCCCCBBBAAAA99999988899AAA99888888889888999888888999A99A988788777788888888999999A99AAA999888778888899AA989887777765545443222022222222222222222222222000000000000000000000000000000000000000000000000000000000000002222222453222222222233444555555565678ABBCCCCCECECCECECCCBA987554222222222222232222322222222222222222222222222222222232223223223232232222222222222220222222049B989888888888777885445555555447BEECB842233222220000220000002555445754345554357ACAA87322222222222222222222222EECEECCCCCCCCCBBBAAAA99999988899AAA99888888889888999888888999A99A988788777788888888999999A99AAA999888778888899AA989887777765545443222022222222222222222222222000000000000000000000000000000000000000000000000000000000000002222222453222222222233444555555565678ABBCCCCCECECCECECCCBA987554222222222222232222322222222222222222222222222222222232223223223232232222222222222220222222049B989888888888777885445555555447BEECB842233222220000220000002555445754345554357ACAA87322222222222222222222222;
		rom_data[39] <= 3840'hCCCCCCCBBBBAA998888888899A999998888899999999888888989999988888887777888889998999A999AAA99988777888889AA9999888877777655544322220202202022022222222232223220000000000000000000000000000000000000000000000000000000020000002220000200022223344444555555577889BCCCCBBBCCCCBAAACC9889A864322222222222222222232222222222222222222222222322232222223223222232222222222202202222220238BA89998887888888885444555555457CEECBA86532222000022232200000355434443220222222247989A600322222222222222222222EEECCECCCCCCCCCBBBBAA998888888899A999998888899999999888888989999988888887777888889998999A999AAA99988777888889AA9999888877777655544322220202202022022222222232223220000000000000000000000000000000000000000000000000000000020000002220000200022223344444555555577889BCCCCBBBCCCCBAAACC9889A864322222222222222222232222222222222222222222222322232222223223222232222222222202202222220238BA89998887888888885444555555457CEECBA86532222000022232200000355434443220222222247989A600322222222222222222222;
		rom_data[40] <= 3840'hBCBCCCCBBAAAA9998888888888999999888888999A99888888888998888888887777888888998999A999AAA99998877777899A9A99888887778887775533222222222220222022222232233232000000000000000002020000000000000000000000000000000000020000000200000000000222233333345555555778899BCCBBCCCBB9888AB6578ACB987532222222222322222222222222220220222222222222222323232222232322223222222222222222222227EEA9898888888878896444454555445CEEEC98887335643334457753300224433444322222333322027789620222222222222222222222EECCCBBBBCBCCCCBBAAAA9998888888888999999888888999A99888888888998888888887777888888998999A999AAA99998877777899A9A99888887778887775533222222222220222022222232233232000000000000000002020000000000000000000000000000000000020000000200000000000222233333345555555778899BCCBBCCCBB9888AB6578ACB987532222222222322222222222222220220222222222222222323232222232322223222222222222222222227EEA9898888888878896444454555445CEEEC98887335643334457753300224433444322222333322027789620222222222222222222222;
		rom_data[41] <= 3840'hBBBBCBCBAAA99A999988888888889999888889999A9988888888898888889888878888888999999AA999AABBAA98877777889BA999888887678889986533320202022222222222222222322332200000222333322233333222200000000000000000000000000000000000000000000000002022222333443444455788889AAA9ABBABB98766545678ACCCEB9775432222222232222222222222222222222222222232222222232322223222222222222222222202025CEC98888888889877875434445444458EEEEA8899536AA87778888888755554222334333234543344223899830322222222222222222222CCBCBBBBBBBBCBCBAAA99A999988888888889999888889999A9988888888898888889888878888888999999AA999AABBAA98877777889BA999888887678889986533320202022222222222222222322332200000222333322233333222200000000000000000000000000000000000000000000000002022222333443444455788889AAA9ABBABB98766545678ACCCEB9775432222222232222222222222222222222222222232222222232322223222222222222222222202025CEC98888888889877875434445444458EEEEA8899536AA87778888888755554222334333234543344223899830322222222222222222222;
		rom_data[42] <= 3840'hBBBBBBBAAA999AAAA99998888888899888788999999988878888899888888888778888888999989999999ABBBA99887777899ABA9988887667888898753333222222202020202222222232323322002223333332233333333332220000000000000000020000000000000000000000000000200202222323333434579A998A9889A9ABBA87554577778999ABCCCC987533222222232222222222222222222222232222323232322232322323222222222222202222227EC98889988899877764334444444448CECBA889A86678766777777788888753222022323343333323544588B73222222222222222222222BBBBBBBBBBBBBBBAAA999AAAA99998888888899888788999999988878888899888888888778888888999989999999ABBBA99887777899ABA9988887667888898753333222222202020202222222232323322002223333332233333333332220000000000000000020000000000000000000000000000200202222323333434579A998A9889A9ABBA87554577778999ABCCCC987533222222232222222222222222222222232222323232322232322323222222222222202222227EC98889988899877764334444444448CECBA889A86678766777777788888753222022323343333323544588B73222222222222222222222;
		rom_data[43] <= 3840'hBBBBAAAAAAA9A9A999A998888888788888788888999888777888898888788888777778888999999999989AABBA99999887889AB99888876578898888753444322022222222222222223223233222022233332333333333333333332220000000000000000200000000000000000000000000000020222222233334589998788889888888755567787887789999BBBBCC9743222222222222222222222222222222232322222222322222322223222222222222222223AC97788888899877754334444444436BEA888898755656566777778787888742220002223433232323345434884222222222222222222222CBBBBABBBBBBAAAAAAA9A9A999A998888888788888788888999888777888898888788888777778888999999999989AABBA99999887889AB99888876578898888753444322022222222222222223223233222022233332333333333333333332220000000000000000200000000000000000000000000000020222222233334589998788889888888755567787887789999BBBBCC9743222222222222222222222222222222232322222222322222322223222222222222222223AC97788888899877754334444444436BEA888898755656566777778787888742220002223433232323345434884222222222222222222222;
		rom_data[44] <= 3840'h9AAAA99999A999A9A99998888888777877788888898877778888988888888888777778888889A999898889ABA9999AA9878889A98888865578998788754454422222022022022022222232323322223333233232323232333233333323202000000000000220000000000002220000000000000002022022234445678877677787756565555567777754468888889ABCECA9753222222222222222222222222222222232323232223232222322222222222022222037CB87788889888777633333333444447AA8788875555556677777888888888620233222223200222022222233454222222222222222222222CCBAA9AA9AAAA99999A999A9A99998888888777877788888898877778888988888888888777778888889A999898889ABA9999AA9878889A98888865578998788754454422222022022022022222232323322223333233232323232333233333323202000000000000220000000000002220000000000000002022022234445678877677787756565555567777754468888889ABCECA9753222222222222222222222222222222232323232223232222322222222222022222037CB87788889888777633333333444447AA8788875555556677777888888888620233222223200222022222233454222222222222222222222;
		rom_data[45] <= 3840'h88899899999999999988888888877777778878888888777788998988888888887757788888899A98888889A988899AA987889A99888886557999888885555453222222222022222222232323233333333233233333333332333323333232222220000000000000000000000020000000000000000022020223345655557777787554576555445566754334788878889ABCCECCB974322022222222222222222322323222323232322222323222322222222222222238CA88878888765665333233444334445775777655555556777888888888888523332433322443000020002244333222222222222222222222ECBBA98888899899999999999988888888877777778878888888777788998988888888887757788888899A98888889A988899AA987889A99888886557999888885555453222222222022222222232323233333333233233333333332333323333232222220000000000000000000000020000000000000000022020223345655557777787554576555445566754334788878889ABCCECCB974322022222222222222222322323222323232322222323222322222222222222238CA88878888765665333233444334445775777655555556777888888888888523332433322443000020002244333222222222222222222222;
		rom_data[46] <= 3840'h78888888888898998888888888877777777878888888888888999988898988988777788878899998878889987789AA998888999888888655899998898655555432220220222222222222223233233332333333323232323333333323232323222220000000000000000000000000000000000000000020222222455555677677764348544553455555534456777788889AABCEEECA975442222222222222222222222323222322323232322232222222222222222239C988766777665543223333333344444455555555555677788888888989888532345544565798567432202244354222223222232222222222BCBBA98878888888888898998888888888877777777878888888888888999988898988988777788878899998878889987789AA998888999888888655899998898655555432220220222222222222223233233332333333323232323333333323232323222220000000000000000000000000000000000000000020222222455555677677764348544553455555534456777788889AABCEEECA975442222222222222222222222323222322323232322232222222222222222239C988766777665543223333333344444455555555555677788888888989888532345544565798567432202244354222223222232222222222;
		rom_data[47] <= 3840'h88887777878888888888878888777777777887878788888888999989889988988887888778899888878889877789AA9A988898888888765789AA999986555555432222022220222222232323233323233232323323333332332333333232222222222000000000000000000000000000000000000000000220203334554555555542343344444455555555556777777788888ACCCCEECBA8754222222222222223232232232232322222232222222222222222202027A9877677766543222232333334444454445555555567788888999999999973223454557889888AC766543222454222222223222222222232BBBBAA9988887777878888888888878888777777777887878788888888999989889988988887888778899888878889877789AA9A988898888888765789AA999986555555432222022220222222232323233323233232323323333332332333333232222222222000000000000000000000000000000000000000000220203334554555555542343344444455555555556777777788888ACCCCEECBA8754222222222222223232232232232322222232222222222222222202027A9877677766543222232333334444454445555555567788888999999999973223454557889888AC766543222454222222223222222222232;
		rom_data[48] <= 3840'h8888877777777778888887787777777777777777778888888899999899988889888888888898988888888888888AAA9AA98888888887766788AAAAA976565556654322222222202222222223232333323233323232323233233332333232322222222200000000000000000000000000000000000020220020020022333455555433002334444454455566556667776677777898899BCCEEECA865432222222222222322323223232323223232232222222222222224798899887553322222233333334444444455555556778889999A9AAAAAAA844445555677787578888BB96220233222322222222222322222ABBBBB998888877777777778888887787777777777777777778888888899999899988889888888888898988888888888888AAA9AA98888888887766788AAAAA976565556654322222222202222222223232333323233323232323233233332333232322222222200000000000000000000000000000000000020220020020022333455555433002334444454455566556667776677777898899BCCEEECA865432222222222222322323223232323223232232222222222222224798899887553322222233333334444444455555556778889999A9AAAAAAA844445555677787578888BB96220233222322222222222322222;
		rom_data[49] <= 3840'h99998877777767787788877787777777778777777778878888898989999988888888888888998888888889998889A9999987887787777767789BBB997777777887652222022222222223232323232323332323232323323233233332323222222222222200000000000000000000000000000000002220202000000022233445433322223434333445455555556666556776777788899AABCCEECBB98532222222223222232323223232322222222222222222222222588AA975432222222323233334444454555555556778889AAABABAAAABBB8577677787888767775578998532022223222322222223222322AABBBA9999998877777767787788877787777777778777777778878888898989999988888888888888998888888889998889A9999987887787777767789BBB997777777887652222022222222223232323232323332323232323323233233332323222222222222200000000000000000000000000000000002220202000000022233445433322223434333445455555556666556776777788899AABCCEECBB98532222222223222232323223232322222222222222222222222588AA975432222222323233334444454555555556778889AAABABAAAABBB8577677787888767775578998532022223222322222223222322;
		rom_data[50] <= 3840'h999888887777778878887877777777778778777777777788888888899A998788888887788899888899989999998999999987777776667777679BBA99889888998875422222220222222222323333233323323232323233333332323333232322222222222200000000000000000000000000000000222220020000000000223333322222333332234454445555555555667676667788899A999BBCCEEEA87655432222222223223222232323232232222222222222223556542222222222223233333334444455555556778889AABBBBBBBCBBB844577657778888766422323477897322222222222232222222229AAAA998999888887777778878887877777777778778777777777788888888899A998788888887788899888899989999998999999987777776667777679BBA99889888998875422222220222222222323333233323323232323233333332323333232322222222222200000000000000000000000000000000222220020000000000223333322222333332234454445555555555667676667788899A999BBCCEEEA87655432222222223223222232323232232222222222222223556542222222222223233333334444455555556778889AABBBBBBBCBBB84457765777888876642232347789732222222222223222222222;
		rom_data[51] <= 3840'h88877778777878888777778877777888887777877778778888888888998988787877777788989888989999A9998899999998877776667777789AA88999999AA98875432220222222222232323232332332322323232332323233333232232222222222222222200000000000000000000000000000202002000000000002222222222222323332223344444455555555556555656677889888899998ABCCCCCBB965567533322222232222322223222222222222220222222222222222222223323334444455555555667888AAABBBCCCCCCCA524555767877887787400000000226BC52222232322322223223229998888888877778777878888777778877777888887777877778778888888888998988787877777788989888989999A9998899999998877776667777789AA88999999AA98875432220222222222232323232332332322323232332323233333232232222222222222222200000000000000000000000000000202002000000000002222222222222323332223344444455555555556555656677889888899998ABCCCCCBB965567533322222232222322223222222222222220222222222222222222223323334444455555555667888AAABBBCCCCCCCA524555767877887787400000000226BC5222223232232222322322;
		rom_data[52] <= 3840'h877667777777778888887878877788888777888777887788888888898988888888887777888888888999A9AA99999AAA9898877776667777789A98899999BBB99865542222202222222222232323232323232323232323323323232323322222222222202222222220202222022000000000000000200200200000000000000000202022223333333333334445445555555555567667777777777888899999ABCBA9AACCB9985555332222222222222222222222222222220222222222222232233333344444555555678899AABBCCCCCCCEB533555567864553335543000000000049B752323223222322232232AA987888877667777777778888887878877788888777888777887788888888898988888888887777888888888999A9AA99999AAA9898877776667777789A98899999BBB99865542222202222222222232323232323232323232323323323232323322222222222202222222220202222022000000000000000200200200000000000000000202022223333333333334445445555555555567667777777777888899999ABCBA9AACCB9985555332222222222222222222222222222220222222222222232233333344444555555678899AABBCCCCCCCEB533555567864553335543000000000049B752323223222322232232;
		rom_data[53] <= 3840'h8756677777777777887788888777889888888888788888888888889898888888888887778888888889999AAA9889AABA988887777677775678AAAAAA9999ABA998755432222222022222323232323232323232323232323323233232322322222222222222220222022220222222222020000000000000020000000000000002200002020222222233333433444555555555555566666665576777778888888899999ABCCCCCAABB86665443322222220200200002020202220222222222222222233344445555555677899AABCCCCEEECA974345555544220220020200000022200026996323322232223222322AA9878888756677777777777887788888777889888888888788888888888889898888888888887778888888889999AAA9889AABA988887777677775678AAAAAA9999ABA998755432222222022222323232323232323232323232323323233232322322222222222222220222022220222222222020000000000000020000000000000002200002020222222233333433444555555555555566666665576777778888888899999ABCCCCCAABB86665443322222220200200002020202220222222222222222233344445555555677899AABCCCCEEECA974345555544220220020200000022200026996323322232223222322;
		rom_data[54] <= 3840'h7656777767777777777888888888899988889988888887788878889999888888888888788888888889999A998989ABBCA98888767777666689ABBBBBA999A9A9A98655432220222222222232323232323232232223222323232323323232322222222222202222222220222202022222222000000000000000000000000000020202000200022022222333333444444554444455556555555666666677878877888888ABCCBABBCCBBCCBA988877676554543444445555555554333344554444434444334445555677889AABCCCEEECA975554434444320000020022000002220202202489754332223232232232999877877656777767777777777888888888899988889988888887788878889999888888888888788888888889999A998989ABBCA98888767777666689ABBBBBA999A9A9A98655432220222222222232323232323232232223222323232323323232322222222222202222222220222202022222222000000000000000000000000000020202000200022022222333333444444554444455556555555666666677878877888888ABCCBABBCCBBCCBA988877676554543444445555555554333344554444434444334445555677889AABCCCEEECA975554434444320000020022000002220202202489754332223232232232;
		rom_data[55] <= 3840'h666667677767777777888888988899988899999888887777888889999999888888888888888888888899A998888AABCCB9889877778766778AABBCCBA9A9999ABBA8777422222222222232232323232323223223222322323232332323232222222222222222220220222202222202220222220000000000000000000000000202200000000000000022222223343444544344445555555565655556567777778888889999899A99ABC99999CCCAAABB99AA9A89A98888787875554455677788889985666555545667777777889988654344444344343000000022422220233320025522369A832222222322322288887777666667677767777777888888988899988899999888887777888889999999888888888888888888888899A998888AABCCB9889877778766778AABBCCBA9A9999ABBA8777422222222222232232323232323223223222322323232332323232222222222222222220220222202222202220222220000000000000000000000000202200000000000000022222223343444544344445555555565655556567777778888889999899A99ABC99999CCCAAABB99AA9A89A98888787875554455677788889985666555545667777777889988654344444344343000000022422220233320025522369A8322222223223222;
		rom_data[56] <= 3840'h555555556666777778888888989899988899AA998888777777888888888888888888888788899998888998888899ABCBBA988887778777788ABAABBBAABAA99BCCCBA9973222202222222232232323232232222223223223233232332322322222222222222222222222022220222222222222222200000000000000000000002020000000000000000002022232333444444433455565555555555556666678878888887788888888866777899999A99ACCB99899777778755445545557889ABCCB878887754445555554444555422333444443444520000000244443454554430037522358953232232232223277887665555555556666777778888888989899988899AA998888777777888888888888888888888788899998888998888899ABCBBA988887778777788ABAABBBAABAA99BCCCBA9973222202222222232232323232232222223223223233232332322322222222222222222222222022220222222222222222200000000000000000000002020000000000000000002022232333444444433455565555555555556666678878888887788888888866777899999A99ACCB99899777778755445545557889ABCCB8788877544455555544445554223334444434445200000002444434545544300375223589532322322322232;
		rom_data[57] <= 3840'h5555554555676767888889898898998888899A9987777777778888877788888888889887888999888888888888889AAAA9988887788777889AAAAABBBBBAA9ACCECCBBB85320222222223223232323232322322222222323232332323232222222222222222220220222220222220222222222222222200000000000000000000002000000000000000000020222332333344343554555555555555555555677767777766665676777777776567889866787654556566777543335566556777989985687755555445554444444554334554445544444220022223344445545445553024333337A74322222223223877776555555554555676767888889898898998888899A9987777777778888877788888888889887888999888888888888889AAAA9988887788777889AAAAABBBBBAA9ACCECCBBB85320222222223223232323232322322222222323232332323232222222222222222220220222220222220222222222222222200000000000000000000002000000000000000000020222332333344343554555555555555555555677767777766665676777777776567889866787654556566777543335566556777989985687755555445554444444554334554445544444220022223344445545445553024333337A74322222223223;
		rom_data[58] <= 3840'h444544445566667778888888998989988889AA988877777777888887777888878888888778899988888888888887899889988777888778888899AABBBBBA99ACCEECCCBA84222222222222232323232322322232232322232232323232223222222222222222222222020222022222220222222222222222200000000000000000000000000000000000000202222322222334445555555555555445555555655555565555555555677667755577777555555555555577654434445666777778988878765555554455543344344554455555545555434433554454222345444455663233356358AA75333232222287775555444544445566667778888888998989988889AA988877777777888887777888878888888778899988888888888887899889988777888778888899AABBBBBA99ACCEECCCBA84222222222222232323232322322232232322232232323232223222222222222222222222020222022222220222222222222222200000000000000000000000000000000000000202222322222334445555555555555445555555655555565555555555677667755577777555555555555577654434445666777778988878765555554455543344344554455555545555434433554454222345444455663233356358AA753332322222;
		rom_data[59] <= 3840'h54454455556666677888888888989988888999888777787877888877788877778888988778899988898888888877788878887777787778888889BBAAABBA9AABCCECCBBB9532222222222323232323223222322222222322323232323232222222222222220222222222222222202222222222222222222222220000000000000000200000000000000000000202222222222334455555444555544545455545445455555555555555556885456677655555565556657754444445566776777898998755555544586653222344455444555544455530584443454300022333345555544334854578A988764455328775555554454455556666677888888888989988888999888777787877888877788877778888988778899988898888888877788878887777787778888889BBAAABBA9AABCCECCBBB9532222222222323232323223222322222222322323232323232222222222222220222222222222222202222222222222222222222220000000000000000200000000000000000000202222222222334455555444555544545455545445455555555555555556885456677655555565556657754444445566776777898998755555544586653222344455444555544455530584443454300022333345555544334854578A98876445532;
		rom_data[60] <= 3840'h55554445566667777788888888888988999887777788888877788888888877777788898888899989998899998877788887777777778788887789AB9ABBCAAAABCCCCCCBAA7322202222222223232323222322222222322223223232232223222222222222222222202222220222222222222222222222222222222220000000000000000000000000000000000220020222223323335544344455454454555444454455555555544444467645666555555555555655665545554565456556679888876655544333544322224554444544355444555302334555554320002322344455554346445789A9879BCB8528876555555554445566667777788888888888988999887777788888877788888888877777788898888899989998899998877788887777777778788887789AB9ABBCAAAABCCCCCCBAA7322202222222223232323222322222222322223223232232223222222222222222222202222220222222222222222222222222222222220000000000000000000000000000000000220020222223323335544344455454454555444454455555555544444467645666555555555555655665545554565456556679888876655544333544322224554444544355444555302334555554320002322344455554346445789A9879BCB852;
		rom_data[61] <= 3840'h55544444555666677778888888888888888877777788888887888888888877778778888888989999999999A98775678887777777777888887789A999BCCBBAAABCECCCBAA8532022222222322323232323222222222222322323223232322222222222222222222222022022220220220222222222222222222222222200000000000000000000000000000000000000202222222234544433355544444555554454555555555555444420345555555455555545555556555555554455555688888765555543247543322234545444443455545555420235555555432034443355555554447435678875568879CA8887656555544444555666677778888888888888888877777788888887888888888877778778888888989999999999A98775678887777777777888887789A999BCCBBAAABCECCCBAA8532022222222322323232323222222222222322323223232322222222222222222222222022022220220220222222222222222222222222200000000000000000000000000000000000000202222222234544433355544444555554454555555555555444420345555555455555545555556555555554455555688888765555543247543322234545444443455545555420235555555432034443355555554447435678875568879CA;
		rom_data[62] <= 3840'h55555444445555556677777777778877877788877788888888899A998887778887777888899989999889AAAA88555578877877788778888767889899ACCCBAAABBCCCCBA99742222222222232322322322232222222222232232232232223222222222222222202222222222222222222222222222222222222222222222202000000000000000000000000000000000000222222223233433345533344455454445555455554454444332345554544454554434545555555555554555455788887665555433335333323443544444444434544555422235567544443345555445664554445555777777577899998888766555555444445555556677777777778877877788877788888888899A998887778887777888899989999889AAAA88555578877877788778888767889899ACCCBAAABBCCCCBA9974222222222223232232232223222222222223223223223222322222222222222220222222222222222222222222222222222222222222222220200000000000000000000000000000000000022222222323343334553334445545444555545555445444433234555454445455443454555555555555455545578888766555543333533332344354444444443454455542223556754444334555544566455444555577777757789999;
		rom_data[63] <= 3840'h545544444444555555566777777777777878888888888888999AAA999887778887767778898888998899AAAA98644578888888888777887656778889ACCCBBAABBBBCCCBBA9742222222223222323232222222222232222223223223223222222222222222222222202222022220222222222222222222222222222222222222220000000000000000000000000000000002222222220233323333334433343444455544455544444444434444444444444442245555555555555455544467788765555554343202444445444444333444455555545354225555444334576543348634433335667777679A66887687887755545544444444555555566777777777777878888888888888999AAA999887778887767778898888998899AAAA98644578888888888777887656778889ACCCBBAABBBBCCCBBA9742222222223222323232222222222232222223223223223222222222222222222222202222022220222222222222222222222222222222222222220000000000000000000000000000000002222222220233323333334433343444455544455544444444434444444444444442245555555555555455544467788765555554343202444445444444333444455555545354225555444334576543348634433335667777679A668876;
		rom_data[64] <= 3840'h4444544444444555455566677777777788888888888998899A99AA99888778888777778988888899889AAAA998754577877788889877776567678889BCCBBBAABAABBBCCCBCA732222222222323223222232222222222222222223223223232222222222222222222220222220222222222222222222222222222222222222222222200000000000000000000000000000000222220202232222333333332333345544434434344432454433333355554454323345554445455554433344567778754665544530233454454544434444445565445444430043344343334554442343333223346677755577557865888876544444544444444555455566677777777788888888888998899A99AA99888778888777778988888899889AAAA998754577877788889877776567678889BCCBBBAABAABBBCCCBCA732222222222323223222232222222222222222223223223232222222222222222222220222220222222222222222222222222222222222222222222200000000000000000000000000000000222220202232222333333332333345544434434344432454433333355554454323345554445455554433344567778754665544530233454454544434444445565445444430043344343334554442343333223346677755577557865;
		rom_data[65] <= 3840'h444444455555555555567777777777788888999899A999899A999888888888888878788988778898889AAA988876555665557888897777777767888ABCBBBABBBABBAABBCCCC95222222232322322223222222222222222323223223232322222222222222222222022222202222022222222222223222222222322222222220222222220000000000000000000000000000000222220222220333322233222245543233233344432234333322234544434432334444333445544533334456777875566554554333335445443334445545555554555432024023433233334444300222202355556655342456765788887544444444455555555555567777777777788888999899A999899A999888888888888878788988778898889AAA988876555665557888897777777767888ABCBBBABBBABBAABBCCCC952222222323223222232222222222222223232232232323222222222222222222220222222022220222222222222232222222223222222222202222222200000000000000000000000000000002222202222203333222332222455432332333444322343333222345444344323344443334455445333344567778755665545543333354454433344455455555545554320240234332333344443002222023555566553424567657;
		rom_data[66] <= 3840'h3344444445555555566777787877877888899A99AAAA99899999888888889988888877899877789888899998888765555545678889887777876689AAABBBAAAABBAAA9AAABCCC82222222222322323223222222222222222222223232322223222222222222222222222222222222202222222222222222223222222222222222022022222220000000000000000000000020200223200220223333223232222454322222223433202222222222333333333333334344333444334333553477678755553443333434355543223444543332234544553232230033333334343202023300345655565544344575557888886543344444445555555566777787877877888899A99AAAA99899999888888889988888877899877789888899998888765555545678889887777876689AAABBBAAAABBAAA9AAABCCC82222222222322323223222222222222222222223232322223222222222222222222222222222222202222222222222222223222222222222222022022222220000000000000000000000020200223200220223333223232222454322222223433202222222222333333333333334344333444334333553477678755553443333434355543223444543332234544553232230033333334343202023300345655565544344575557;
		rom_data[67] <= 3840'h4344444455555556677777888878888888889AAAABAAA999AA98888888899999988887889887788887889998788765455544567789987787777789AAAABBAAA9A99AA999AACEE94222222222223222222222222222222222322323222223222222222222222222222022202222222222222222222222322322222222222222222222222222222222000000000000000000000002022202222222222222222002332220222233233220000222020222222323222233334433333333333542345665544433433233333234433233345420000000333454333320023334455422202233002344445555555565555556888887654344444455555556677777888878888888889AAAABAAA999AA98888888899999988887889887788887889998788765455544567789987787777789AAAABBAAA9A99AA999AACEE94222222222223222222222222222222222322323222223222222222222222222222022202222222222222222222222322322222222222222222222222222222222000000000000000000000002022202222222222222222002332220222233233220000222020222222323222233334433333333333542345665544433433233333234433233345420000000333454333320023334455422202233002344445555555565555556;
		rom_data[68] <= 3840'h44454444445556567777788888888988889899AABBAAAA9A9999988889899AA9999988888888888877778887788755455555677788887777777889AAAABBBBA99999A9989ACCEB62222222223223232322222222222222222222232323223222322222222222222222222222202222222222222223222222222232222222222222222220222222222220000000000000000000002202222322222222022220200002020022222223220000020220200222222233333333333223322223323456545533343222022320223333333432000000000233343552022232233432222002200222344345555555576554558888887544454444445556567777788888888988889899AABBAAAA9A9999988889899AA9999988888888888877778887788755455555677788887777777889AAAABBBBA99999A9989ACCEB6222222222322323232222222222222222222223232322322232222222222222222222222220222222222222222322222222223222222222222222222022222222222000000000000000000000220222232222222202222020000202002222222322000002022020022222223333333333322332222332345654553334322202232022333333343200000000023334355202223223343222200220022234434555555557655455;
		rom_data[69] <= 3840'h54454445545555556777788888899998889999AABAAAAAAAA99888999999AAAA999888888988888887778876577655445567777778887777778889A9AABCCBA9999999888ACEEC84222222222232222222222222222222222222322322322232222222222222222222222222222222222222222222222232232222222222222222022222222222222222222000000000000000202020222202022220022000000022200202200002000002020020002022022223223323222222222333223456555534332222022220222223334320000000000002223453000243322022220000000222433575455555556543338888888754454445545555556777788888899998889999AABAAAAAAAA99888999999AAAA999888888988888887778876577655445567777778887777778889A9AABCCBA9999999888ACEEC8422222222223222222222222222222222222232232232223222222222222222222222222222222222222222222222223223222222222222222202222222222222222222200000000000000020202022220202222002200000002220020220000200000202002000202202222322332322222222233322345655553433222202222022222333432000000000000222345300024332202222000000022243357545555555654333;
		rom_data[70] <= 3840'h7555444555555555677778888899999989999AAA9AAAAABB99899999A9AAABAAA9988888989888998767787655655554557888887788877788899889ABBCCBB9888888889ACCECB522222222222222222222222222222222222223223223222222322222222222222222222222222222222222232223222322232222322222222222220222222222223232222000000000000000220222200000000000020000200000000000000000000000200200000222022222220222020200322322355555433222222220222022002334320000000000000022223320002330000023200000222332355434555555553022888888887555444555555555677778888899999989999AAA9AAAAABB99899999A9AAABAAA9988888989888998767787655655554557888887788877788899889ABBCCBB9888888889ACCECB522222222222222222222222222222222222223223223222222322222222222222222222222222222222222232223222322232222322222222222220222222222223232222000000000000000220222200000000000020000200000000000000000000000200200000222022222220222020200322322355555433222222220222022002334320000000000000022223320002330000023200000222332355434555555553022;
		rom_data[71] <= 3840'h7655445555555556777777787888998988999AAA999AAABB99999999A99AAAABBA988888999888888666787776556665567899887678887778988878ABCCCCBA888877889BCCCCC732222222232223222232222222222222232222322232222222222222222222222222222222022222222222222322222222222223222222222222022222222222222232332222000000000202022200000000000000000000000000000000000000000000002000002000202222202000000000222022333343220220233000020000202354200000000000000002000253000002220220000002233332202344555554543222888888887655445555555556777777787888998988999AAA999AAABB99999999A99AAAABBA988888999888888666787776556665567899887678887778988878ABCCCCBA888877889BCCCCC732222222232223222232222222222222232222322232222222222222222222222222222222022222222222222322222222222223222222222222022222222222222232332222000000000202022200000000000000000000000000000000000000000000002000002000202222202000000000222022333343220220233000020000202354200000000000000002000253000002220220000002233332202344555554543222;
		rom_data[72] <= 3840'h8765555555555556777777778888889888999AA999999ABAA99AA9999A9999ABBB998889999888888766777777767777777889887667888778887668ACCBCCBA99987778ABCCCCB842222222222222222222222222222222222223223222232232223222222222222222222222222222222232232222223232322322222222222222222222222222223223223323200000000002202202000000000000000000000000000000000000000000000000000000000000000002000000000002022222000020222000000000022342000002000000000000000035400000000000000022332232202354575555544233888888888765555555555556777777778888889888999AA999999ABAA99AA9999A9999ABBB998889999888888766777777767777777889887667888778887668ACCBCCBA99987778ABCCCCB842222222222222222222222222222222222223223222232232223222222222222222222222222222222232232222223232322322222222222222222222222222223223223323200000000002202202000000000000000000000000000000000000000000000000000000000000000002000000000002022222000020222000000000022342000002000000000000000035400000000000000022332232202354575555544233;
		rom_data[73] <= 3840'h8876656555556557787777777888899888899AA99999999A99ABA9999999889AAAA999AAA999988887777776777888887778889877679988777775579BBBCCCBAAA987789BBBCCBA63222222222322232222222222222222222322232232322222222222222222222222222222222222222222322323232222223222222222222222222222222222322232232323332000000222322200000000000000000000000000000000000000000000000000000000000000000000000000000000000020000200000000000000020220000022022222000000000002520000000000000022322222333322357555554333888888888876656555556557787777777888899888899AA99999999A99ABA9999999889AAAA999AAA999988887777776777888887778889877679988777775579BBBCCCBAAA987789BBBCCBA63222222222322232222222222222222222322232232322222222222222222222222222222222222222222322323232222223222222222222222222222222222322232232323332000000222322200000000000000000000000000000000000000000000000000000000000000000000000000000000000020000200000000000000020220000022022222000000000002520000000000000022322222333322357555554333;
		rom_data[74] <= 3840'h88887765555666677778777778889888888889A99999888A9AAAA9999999888899999BCCBAA99887777777766778888888878889877899887776555689ABCCCCBBAA88789AAABBBB842222222222222222222222222222222222322232222222223222222322222222222222222222222222222322222222323222223222222222222222222222222232323232323232000022323322000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002233202020000000000000000000000000022222223300000246555553238888888888887765555666677778777778889888888889A99999888A9AAAA9999999888899999BCCBAA99887777777766778888888878889877899887776555689ABCCCCBBAA88789AAABBBB84222222222222222222222222222222222232223222222222322222232222222222222222222222222222232222222232322222322222222222222222222222223232323232323200002232332200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000223320202000000000000000000000000002222222330000024655555323;
		rom_data[75] <= 3840'h88888775555666777777777778898888888888999988888999999999889988778899ABCCBA9887777777788877778888888777898887898866665455889BBCCCBBA99888899AABBBA52222222322232222222222222222222222222222323223222223222222222222222222222222222223232223232323222232232222222222222222222222323223232323233232222232222320020000002200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000002002020200200000000000000000000002320222220000000002555554338888888888888775555666777777777778898888888888999988888999999999889988778899ABCCBA9887777777788877778888888777898887898866665455889BBCCCBBA99888899AABBBA5222222232223222222222222222222222222222232322322222322222222222222222222222222222323222323232322223223222222222222222222222232322323232323323222223222232002000000220000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000200202020020000000000000000000000232022222000000000255555433;
		rom_data[76] <= 3840'h888888755555677777777767788988888888889988888888998999988888888778889BBA988887777777788988766788888766899988888755555445789ABCCBAA888887799AAAABA742222222222222222222222222222222232232322223222222223232223222222222222222222223222232323232223232232222322222222222222222222223232232323323333222322002200020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000245220000000000000002344432388888888888888755555677777777767788988888888889988888888998999988888888778889BBA988887777777788988766788888766899988888755555445789ABCCBAA888887799AAAABA7422222222222222222222222222222222322323222232222222232322232222222222222222222232222323232322232322322223222222222222222222222232322323233233332223220022000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000002452200000000000000023444323;
		rom_data[77] <= 3840'h888888766766677777776767788888888888889888888888888898887778877777888988888888888788788888767777788776789888888755555544688ABCCA98888977788AAA9A98522222222222222222222222222222222222222232222223223222223222222222222222222222222322222322223222223223232222222222222222222223222323232332322222332200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002B8002000000000000000023332288888888888888766766677777776767788888888888889888888888888898887778877777888988888888888788788888767777788776789888888755555544688ABCCA98888977788AAA9A98522222222222222222222222222222222222222232222223223222223222222222222222222222222322222322223222223223232222222222222222222223222323232332322222332200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002B80020000000000000000233322;
		rom_data[78] <= 3840'h8888887777777677777777777887888778778888777888888888888876677777777788888788899988988888887777777778887898889998555554445789BCCB889999877889999998632222222222222222222222222222222322323222323222322232322222322322222322232223232223323232323232322322222322222222222222222322232232323323233220202200000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002640020000000022000000023222888888888888887777777677777777777887888778778888777888888888888876677777777788888788899988988888887777777778887898889998555554445789BCCB889999877889999998632222222222222222222222222222222322323222323222322232322222322322222322232223232223323232323232322322222322222222222222222322232232323323233220202200000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002640020000000022000000023222;
		rom_data[79] <= 3840'h8888888888777777777778888888877777777777777788888777778765566777666788888889AABAAABBA988888778877788888898888998765656555789BCCB999A9A987789999888752222222232222222222222222222232223222232222232223223223232222223232223222232222322232232323232323223232223222222222222232223223232323232345532000000000022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000022200000000222888888888888888888777777777778888888877777777777777788888777778765566777666788888889AABAAABBA988888778877788888898888998765656555789BCCB999A9A987789999888752222222232222222222222222222232223222232222232223223223232222223232223222232222322232232323232323223232223222222222222232223223232323232345532000000000022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000022200000000222;
		rom_data[80] <= 3840'h888887899987888888778888889887777777777788777878888777887678877777778888888ABBCBCBCCCBA8888778888877888888888899877777767789BCBAA99999A8878999887887322222222222222222222222222222232222322232322232323232232232232222222222222223232322322232232232232322232223222222222222222232323233233233785200000200002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022020000000000002089898888888887899987888888778888889887777777777788777878888777887678877777778888888ABBCBCBCCCBA8888778888877888888888899877777767789BCBAA99999A88789998878873222222222222222222222222222222322223222323222323232322322322322222222222222232323223222322322322323222322232222222222222222323232332332337852000002000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000220200000000000020;
		rom_data[81] <= 3840'h888887799988899AA9878888888887777778787888788788888888888788988888888888899AAABBBBAACBA9887778777777776788878888887888877789BBA9899999A9888999887799632222222232222222222222222232232223223222232322323223222322322323232223223232223223223232323232322223222322222222222322323223232332332323574200000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000020200000000000000088998988888887799988899AA9878888888887777778787888788788888888888788988888888888899AAABBBBAACBA9887778777777776788878888887888877789BBA9899999A98889998877996322222222322222222222222222322322232232222323223232232223223223232322232232322232232232323232323222232223222222222223223232232323323323235742000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000202000000000000000;
		rom_data[82] <= 3840'h8888877899988ABCCA88889888888888777778888878878888998888878888888888888899989999A989AA99887887777777766788877778887898877789A998779AA99998888888889A8522222322222222222222222222222223223222323223232232323232222322222223223222222323232322322323223232322322322223223222222232322323232333334532200000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000889898888888877899988ABCCA88889888888888777778888878878888998888878888888888888899989999A989AA99887887777777766788877778887898877789A998779AA99998888888889A8522222322222222222222222222222223223222323223232232323232222322222223223222222323232322322323223232322322322223223222222232322323232333334532200000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000;
		rom_data[83] <= 3840'h8888877789999CEECBA99998888888888877888887877778889888888887778888888889998888888888899888888878877777777777667788789887888899875689999988887778899BA732222222222222222222222222322322232232232322323232323223232223232322222232323232323232323223232323232322222222222222323223232323323323433322200000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000989989888888877789999CEECBA99998888888888877888887877778889888888887778888888889998888888888899888888878877777777777667788789887888899875689999988887778899BA732222222222222222222222222322322232232232322323232323223232223232322222232323232323232323223232323232322222222222222323223232323323323433322200000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		rom_data[84] <= 3840'h88888877789ACCEEECCBAA98899999999888899888877888889888888887778888899999998988888888899988888888888777778776666777788888888889854589A988878777889A9AA8532222222232222222222222222322232223223232323232323232323223222222322323232323232322323232323223232232232323222322322223223232323323233223222200000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008998989888888877789ACCEEECCBAA98899999999888899888877888889888888887778888899999998988888888899988888888888777778776666777788888888889854589A988878777889A9AA853222222223222222222222222232223222322323232323232323232322322222232232323232323232232323232322323223223232322232232222322323232332323322322220000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		rom_data[85] <= 3840'h8888887779BCEEECEEECBA999AABBBAA9A9A99988888888899988899998778888999A9A999998988888999AA9888888988888777888776555667888888888986557999877787778899999853222322222222222222222222222322232323232323232323232323223223232322222323223232323232323232323232322322222223222222232223232323233322222220200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000989999888888887779BCEEECEEECBA999AABBBAA9A9A99988888888899988899998778888999A9A999998988888999AA9888888988888777888776555667888888888986557999877787778899999853222322222222222222222222222322232323232323232323232323223223232322222323223232323232323232323232322322222223222222232223232323233322222220200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		rom_data[86] <= 3840'h888888777ACEEECECEEECBABBBBCCBBBABBAA88998888898999A9999A987788889A9A9999999899889998ABBA98888889888888888777654556898888778998767888875567777888898887322222232222222222222223223222322323232323232323232232323222323223232322323232323232323232323232323232323232222322322323232323232342022233000000000000000000000000000000000000000202020222020222220000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000099999988888888777ACEEECECEEECBABBBBCCBBBABBAA88998888898999A9999A987788889A9A9999999899889998ABBA988888898888888887776545568988887789987678888755677778888988873222222322222222222222232232223223232323232323232322323232223232232323223232323232323232323232323232323232322223223223232323232323420222330000000000000000000000000000000000000002020202220202222200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		rom_data[87] <= 3840'h8888887789CECECEEEEECCCCCCECCCCCCBBB98889988899999A9AA999988789999A9999899999998999899AA9999988889998899888777666777888887889988878876543467778888888874222222222222222222222222322322323232323232323232323232322323223223223232322323233232323233232323232232222223222232232232232323257532223322000000000000000000000000000000333333333333333333333333333322222222323232222220220002020200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000999999988888887789CECECEEEEECCCCCCECCCCCCBBB98889988899999A9AA999988789999A9999899999998999899AA9999988889998899888777666777888887889988878876543467778888888874222222222222222222222222322322323232323232323232323232322323223223223232322323233232323233232323232232222223222232232232232323257532223322000000000000000000000000000000333333333333333333333333333322222222323232222220220002020200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		rom_data[88] <= 3840'h8888887778BCCCEEEEEEEEEEEEEECCCCCCCA98899998999A99A999998988889999999889999999989998888889ACBA9899999999988777777777778888888888877755333357878888887786322322232222222222222222232232232323232323232323232323232323232323232323232323323233323323233232232323232322323223223223232323589543222232000000000000000000000000000003333333433433343333333333333333333333333333333233233323333333222322222223332334455420000222200000000000000000000000000000000000000000000000000000000000000000899998988888887778BCCCEEEEEEEEEEEEEECCCCCCCA98899998999A99A999998988889999999889999999989998888889ACBA9899999999988777777777778888888888877755333357878888887786322322232222222222222222232232232323232323232323232323232323232323232323232323323233323323233232232323232322323223223223232323589543222232000000000000000000000000000003333333433433343333333333333333333333333333333233233323333333222322222223332334455420000222200000000000000000000000000000000000000000000000000000000000000000;
		rom_data[89] <= 3840'h88888877778ACEEEEEEEEECEEEECCECCCCBA99AAAAA999AAA99999888988899A98899999AA9999988988888878ACCA98999A99999888888888777677778888887776433233578877888888885222222222322222223222223223223232323232323232323232323232323223232323232323232332323323323323233232322322232222322322323223578776420002200000000000000000000000000000233333333333333334334334333333333333333333333333333233333323332333333333344555678898854588888773000000000000000000000000000000000000000000000000000000000000009999998988888877778ACEEEEEEEEECEEEECCECCCCBA99AAAAA999AAA99999888988899A98899999AA9999988988888878ACCA98999A9999988888888877767777888888777643323357887788888888522222222232222222322222322322323232323232323232323232323232322323232323232323233232332332332323323232232223222232232232322357877642000220000000000000000000000000000023333333333333333433433433333333333333333333333333323333332333233333333334455567889885458888877300000000000000000000000000000000000000000000000000000000000000;
		rom_data[90] <= 3840'h888888877778ACCEEEEECCEEEEEEECCCBABAA9BBBAAAA9999A9999998898999A9889AAAAAA99898889888888779BA9888899988877888888888788776788888788754333334688778988888973223232222222232222222223223232232323232332332332333233232323232232232323232332323323232332323232323232232232322322232322479B7456420000000000000000000000000000000000333333333333333433333333333333333333333333323232323323232333233333332233334555667888A9AAAAAAABC82000000000000220000000000000000000000000000000000000000000000099899998888888877778ACCEEEEECCEEEEEEECCCBABAA9BBBAAAA9999A9999998898999A9889AAAAAA99898889888888779BA9888899988877888888888788776788888788754333334688778988888973223232222222232222222223223232232323232332332332333233232323232232232323232332323323232332323232323232232232322322232322479B7456420000000000000000000000000000000000333333333333333433333333333333333333333333323232323323232333233333332233334555667888A9AAAAAAABC820000000000002200000000000000000000000000000000000000000000000;
		rom_data[91] <= 3840'h8888887777679ACEECCCCBBCEEEECCCBAAAAAABBBABAA99A99A9999999999899989AAAAAAA998999888999987688888778888777777777788888898766678888887654333335577778998889952222223222222222222232232322323232332332323232332323323232323232323232323232323323333233233323232323223222222232232232237BEB544652000020000000000000000000000000002333333333333434333343343333333333333333323333333333323332332333323332333334455557787888888888889A84200000000038987887677654332220000000000000000000000000000000999989988888887777679ACEECCCCBBCEEEECCCBAAAAAABBBABAA99A99A9999999999899989AAAAAAA998999888999987688888778888777777777788888898766678888887654333335577778998889952222223222222222222232232322323232332332323232332323323232323232323232323232323323333233233323232323223222222232232232237BEB544652000020000000000000000000000000002333333333333434333343343333333333333333323333333333323332332333323332333334455557787888888888889A84200000000038987887677654332220000000000000000000000000000000;
		rom_data[92] <= 3840'h88888877777678ACCBABBBABCCCECCBAABBBBBBBAAAA9999AA9AA998999A9999999A999AA8888998888889887678888877777777776677788888998877767778877775334433467778999888974222322232222223232223222323232323233232332323233233232323223232323223232323232323232332323233233232322322323222323223259CA98544532000000000000000000000000000000233333333333433333343333343343333333333333332333333323332333333333333332323344555677788888888888888A985543202027999AAAABABBAAA987654320000000000000000000000000009998999988888877777678ACCBABBBABCCCECCBAABBBBBBBAAAA9999AA9AA998999A9999999A999AA8888998888889887678888877777777776677788888998877767778877775334433467778999888974222322232222223232223222323232323233232332323233233232323223232323223232323232323232332323233233232322322323222323223259CA98544532000000000000000000000000000000233333333333433333343333343343333333333333332333333323332333333333333332323344555677788888888888888A985543202027999AAAABABBAAA98765432000000000000000000000000000;
		rom_data[93] <= 3840'h8888887777766789999BBAAABCEEECCBBABBBCCBBAA999AAAAAAA998989A99A9889A999A98877888878888887788888776677887777777788888988888877677777787445543357878899877885322222222232232222322232323232323232332323333323323232323232323232323233333333233233232333232332323223222222232232323578B98B83333200000000000000000000000000000233333333333433334333343333333333333333333333333233233323323233233233333333334455567778888888888778878888876553578778788877777766555444333000000000000000000000000999898898888887777766789999BBAAABCEEECCBBABBBCCBBAA999AAAAAAA998989A99A9889A999A98877888878888887788888776677887777777788888988888877677777787445543357878899877885322222222232232222322232323232323232332323333323323232323232323232323233333333233233232333232332323223222222232232323578B98B83333200000000000000000000000000000233333333333433334333343333333333333333333333333233233323323233233233333333334455567778888888888778878888876553578778788877777766555444333000000000000000000000000;
		rom_data[94] <= 3840'h88888887777666777889AAAABCEEEEECBABBBBCBBAAAAAAABAAAA999899999A99999999988777888777788887778887787777777777777888788888778888766666777556754347878888887897322323223222222232223232323232332333323233232332333233232323232323232323232323232332332323333233232322323232322322357998CB78853432020000000000000000000003320233333333333333334333433334343334333333333332333333333233323333333333333323233344555677777777888777777777777677767677777777676655555444332332000000000000000000000009999999888888887777666777889AAAABCEEEEECBABBBBCBBAAAAAAABAAAA999899999A99999999988777888777788887778887787777777777777888788888778888766666777556754347878888887897322323223222222232223232323232332333323233232332333233232323232323232323232323232332332323333233232322323232322322357998CB7885343202000000000000000000000332023333333333333333433343333434333433333333333233333333323332333333333333332323334455567777777788877777777777767776767777777767665555544433233200000000000000000000000;
		rom_data[95] <= 3840'h888888777777666666789ABBBCEEEEECCAAAABBBBBAAAAABABAA9A999989999999999888777777776567887665677778887776767787778887777767888887756566776677755678888788888984222222322322222223232232323233233232333232332332323323323232323232323323233332332333233232323323232232222232322226ABA7589556555432200000000000000000000233333333333333333334333433434433334333333333333333333333333333332333333333333332333455556677777777777777676666555665666666665555555555443433332333200000000000000000000098988888888888777777666666789ABBBCEEEEECCAAAABBBBBAAAAABABAA9A999989999999999888777777776567887665677778887776767787778887777767888887756566776677755678888788888984222222322322222223232232323233233232333232332332323323323232323232323323233332332333233232323323232232222232322226ABA75895565554322000000000000000000002333333333333333333343334334344333343333333333333333333333333333323333333333333323334555566777777777777776766665556656666666655555555554434333323332000000000000000000000;
		rom_data[96] <= 3840'h88888877777666555566789AABCEEEEECA999AABBCBBAAAA9AA9AAAA9998899899889998777877775567875556678777876667777776778877777667787777777767777777777778877778877885322322232223232322232322323323323333323333233233233232332323232323232323323233232323323332332332323222323223222379B95334775687543200000000000000000000033333333333333333343334334334334343333343333333333333333333323323333233333333333333344555666777777777776666555555555556666665555555444434333232322333200000022222222222229999989888888877777666555566789AABCEEEEECA999AABBCBBAAAA9AA9AAAA9998899899889998777877775567875556678777876667777776778877777667787777777767777777777778877778877885322322232223232322232322323323323333323333233233233232332323232323232323323233232323323332332332323222323223222379B9533477568754320000000000000000000003333333333333333334333433433433434333334333333333333333333332332333323333333333333334455566677777777777666655555555555666666555555544443433323232233320000002222222222222;
		rom_data[97] <= 3840'h888888777766655555555778ABCCEEEEBA98999BBBBAA99A99AA9AA9A9989998988888888777777556677755777788776566778888777788877877777767777888877777766788888876788757852232222223222223232323232332332332323323233323323323323332323232323233323323323333323332333233232323232232222358A99533335755855430000000000000000000002233333333333333333333433433434343433343333333333333333333323333333233333333333323333445555666677776666665655555555556656666555544443433333323222232333202223333333333333398989888888888777766655555555778ABCCEEEEBA98999BBBBAA99A99AA9AA9A9989998988888888777777556677755777788776566778888777788877877777767777888877777766788888876788757852232222223222223232323232332332332323323233323323323323332323232323233323323323333323332333233232323232232222358A995333357558554300000000000000000000022333333333333333333334334334343434333433333333333333333333233333332333333333333233334455556666777766666656555555555566566665555444434333333232222323332022233333333333333;
		rom_data[98] <= 3840'h888888777776665555555789ABBBCEECCA98999AAAA99899A9AA9999999899999888887776555665567777567777777765677888887788998888877765556778888877766667887777777875567532232323222323222232232332332332333323323323323323323323233232323232323323323332323332333233323332323232232247AA976433434566533432000000000000000000023333333333333333333433343434343434334333343333333333333333333332333333333333333333333344555556667666665555555555555556666665555443333333232222232222333333333333333323323389989888888888777776665555555789ABBBCEECCA98999AAAA99899A9AA9999999899999888887776555665567777567777777765677888887788998888877765556778888877766667887777777875567532232323222323222232232332332332333323323323323323323323233232323232323323323332323332333233323332323232232247AA9764334345665334320000000000000000000233333333333333333334333434343434343343333433333333333333333333323333333333333333333333445555566676666655555555555555566666655554433333332322222322223333333333333333233233;
		rom_data[99] <= 3840'h8888887777766555555568999BABBCCCCB999899AA9888989A999998988888988888777765555665678877767666677777788888888889999987777765555777777788877667877667777765557532222223222223223232323233333323323233233233233333233233232323323323233233233233333233323332332323232232223578987555444333774224332000000000000000000233333333333333333343334343434343433434343333333333333333333332333323333333333333323334445555565656555555555555555555666666655554333222322222222222323233333333233333332333989888888888887777766555555568999BABBCCCCB999899AA9888989A999998988888988888777765555665678877767666677777788888888889999987777765555777777788877667877667777765557532222223222223223232323233333323323233233233233333233233232323323323233233233233333233323332332323232232223578987555444333774224332000000000000000000233333333333333333343334343434343433434343333333333333333333332333323333333333333323334445555565656555555555555555555666666655554333222322222222222323233333333233333332333;
		rom_data[100] <= 3840'h88888777776666555554577789AABCCCCCA98889999888989999988888887778777776677555677678887766655557887778788888888999A9877776555456666677789877767776677776655576432323232323223222322333232323323333233333233323233233233233332332333233323233323233233332332332333232322357755455544454325853224430000000000000000003333333333333333333334343343433434343434343433333333333333333333333333333333333333333344455555556555555555555555555565666766555443332222222222222222233333333333332332333338988988888888777776666555554577789AABCCCCCA98889999888989999988888887778777776677555677678887766655557887778788888888999A987777655545666667778987776777667777665557643232323232322322232233323232332333323333323332323323323323333233233323332323332323323333233233233323232235775545554445432585322443000000000000000000333333333333333333333434334343343434343434343333333333333333333333333333333333333333334445555555655555555555555555556566676655544333222222222222222223333333333333233233333;
		rom_data[101] <= 3840'h8888777776666555555445455789ABCCCCBA9889AA9A999888999877888766787777777998656776778766777776678877777888889888999877777654455655667777788875566656765675556742323232232223232323232333333323323333233333323333233232332322332332333233233233333233332332332332323223358854334555444433357522332200000000000000000233333333333333333343334343434434343434333333333333333333333333333332333333333333333334345555555555555555555555555565667776655543332222222222222222323333333333333333333333988888888888777776666555555445455789ABCCCCBA9889AA9A999888999877888766787777777998656776778766777776678877777888889888999877777654455655667777788875566656765675556742323232232223232323232333333323323333233333323333233232332322332332333233233233333233332332332332323223358854334555444433357522332200000000000000000233333333333333333343334343434434343434333333333333333333333333333332333333333333333334345555555555555555555555555565667776655543332222222222222222323333333333333333333333;
		rom_data[102] <= 3840'h88887777776655555554444445678ACCCCBA9999BBBBBAA99A9998889988878998877788876666556777788888777888766778998898888988777775334567665667776788766555566656655457532222232223232232323232323233333333233323233323233333333233332332323233233233233233332333332332323323346776543345553333322486300232000000000000000003333333333333333343343433434343443443433434333333333333333333333333333333333333333333344455555555555555555555555556666777776555433222020222022022223233333333333333333333338888888888887777776655555554444445678ACCCCBA9999BBBBBAA99A999888998887899887778887666655677778888877788876677899889888898877777533456766566777678876655556665665545753222223222323223232323232323333333323332323332323333333323333233232323323323323323333233333233232332334677654334555333332248630023200000000000000000333333333333333334334343343434344344343343433333333333333333333333333333333333333333334445555555555555555555555555666677777655543322202022202202222323333333333333333333333;
		rom_data[103] <= 3840'h888777777666655555444443345579BCCCBA888ABCCCBAAAAA99999A99988888988776787766667777888898888888877777888888888788887887754456777655667777787776555556655455575322323223232232323233333333333233233333333333333323323233323233233323323323333333332333333332333322355565333432355322222202453000223000000000000000033333333333343343334334343344344343444343434343333333333333333333333333333333333333333344555555555555545455555555666777777766544333222222222222222223323333333333333333333388988888888777777666655555444443345579BCCCBA888ABCCCBAAAAA99999A999888889887767877666677778888988888888777778888888887888878877544567776556677777877765555566554555753223232232322323232333333333332332333333333333333233232333232332333233233233333333323333333323333223555653334323553222222024530002230000000000000000333333333333433433343343433443443434443434343433333333333333333333333333333333333333333445555555555555454555555556667777777665443332222222222222222233233333333333333333333;
		rom_data[104] <= 3840'h887777777666555555544444333458BCBBBA989ABCCCBBBBAA9AAA9998887787878776777777777877888888888888877778889998888778888887765677777767677677777777765556755555577422322322323223232323232323323333333332333233232333332332333232332332333333323332333332333233232332355533333332244322200020223320023200000000000000233433333333334333333434333434343443434343433333433333333333333333333333333333333333333344455555555555555555555556666777777665544332222222222222222222233333333333333333333388888888887777777666555555544444333458BCBBBA989ABCCCBBBBAA9AAA99988877878787767777777778778888888888888777788899988887788888877656777777676776777777777655567555555774223223223232232323232323233233333333323332332323333323323332323323323333333233323333323332332323323555333333322443222000202233200232000000000000002334333333333343333334343334343434434343434333334333333333333333333333333333333333333333444555555555555555555555566667777776655443322222222222222222222333333333333333333333;
		rom_data[105] <= 3840'h8787777766665555554443433333469BBBCBBAABCBBBBBBCBA9AA999887777777778777788888878888888988888998778888888876567778899887777877787777766677888777776556555555786332323232232323232333323333332332332333233333333233333233233233233233232333333333333333333333332235432233444322333200002000002222020000000000000003433333334333333334333434443444443443434343433433343333333333333333333333333333333333334445555555555555555555555666777777776655443322222222222222222223333334333333333333333888888888787777766665555554443433333469BBBCBBAABCBBBBBBCBA9AA999887777777778777788888878888888988888998778888888876567778899887777877787777766677888777776556555555786332323232232323232333323333332332332333233333333233333233233233233233232333333333333333333333332235432233444322333200002000002222020000000000000003433333334333333334333434443444443443434343433433343333333333333333333333333333333333334445555555555555555555555666777777776655443322222222222222222223333334333333333333333;
		rom_data[106] <= 3840'h88777777766555554544434333333479ABCCCCCCCBCCCBCCBBAAAA999888888777778888889998888888888888889998788888887533456788999887788778888887666788887777665666656556884323232232322323232323333323333333333333333332333233233333233233233233333233333333323333332323233696300234442222222000000200000200000000023000000333333334333333334333434334344343443443444343433343333333333333333333333333333333333333334445555555555555555555556777777777755554333222222222322202232222333333333333333333338888888888777777766555554544434333333479ABCCCCCCCBCCCBCCBBAAAA99988888877777888888999888888888888888999878888888753345678899988778877888888766678888777766566665655688432323223232232323232333332333333333333333333233323323333323323323323333323333333332333333232323369630023444222222200000020000020000000002300000033333333433333333433343433434434344344344434343334333333333333333333333333333333333333333444555555555555555555555677777777775555433322222222232220223222233333333333333333333;
		rom_data[107] <= 3840'h8777777766655555554444333333335789ACCECCCCCCCCECCCAAA9A9A999998887778999998A99877766788888899998877778885322245788998887788878788876655677665666667777665545785322322322323232323333233233323323323323323323333333333233332332332332323333332333333333333233346AC930002232002220000000002000000000000023433333334333343333334334334343434344344343443443443433433343333333333333333333333333434343333334444555555555555555555555667777777666554433222222222222222222222323334333333333333333888888888777777766655555554444333333335789ACCECCCCCCCCECCCAAA9A9A999998887778999998A99877766788888899998877778885322245788998887788878788876655677665666667777665545785322322322323232323333233233323323323323323323333333333233332332332332323333332333333333333233346AC930002232002220000000002000000000000023433333334333343333334334334343434344344343443443443433433343333333333333333333333333434343333334444555555555555555555555667777777666554433222222222222222222222323334333333333333333;
		rom_data[108] <= 3840'h87777777666555555444443433333334578ABCECCCEEECEECBAA9999A9A9A98888888999A88998775544578888899A98877778874302235788887876778888777765555555555567777877755545676543223223223232332323332333333333333333333333333323323323233233233333333333333323333333323334589987420000000000000000000000000000000002333434344333333333343334333434343434344344444444344434344343333333333333333333333333433333343333334444555555555555555555666677777766655543323222222222222222222222333333333333333333338888888887777777666555555444443433333334578ABCECCCEEECEECBAA9999A9A9A98888888999A88998775544578888899A9887777887430223578888787677888877776555555555556777787775554567654322322322323233232333233333333333333333333333332332332323323323333333333333332333333332333458998742000000000000000000000000000000000233343434433333333334333433343434343434434444444434443434434333333333333333333333333343333334333333444455555555555555555566667777776665554332322222222222222222222233333333333333333333;
		rom_data[109] <= 3840'h777777666655555554444333333332333468ABCCCEEECEECCBA99999A9999988888899AA9889887554334789888989988877787642202356777767666778887766555655555555567777776555444578864322323232332332333333233233233233333333333323333332333233233323333333333333333333323335777886443200000000000000000000000000000002334333433333433433433334333434343434443444444444344434434433334343333333333333333333433344343333333434445555555555555555556666777776655554433222222222222222020222233333343333333333333388888887777777666655555554444333333332333468ABCCCEEECEECCBA99999A9999988888899AA98898875543347898889899888777876422023567777676667788877665556555555555677777765554445788643223232323323323333332332332332333333333333233333323332332333233333333333333333333233357778864432000000000000000000000000000000023343334333334334334333343334343434344434444444443444344344333343433333333333333333334333443433333334344455555555555555555566667777766555544332222222222222220202222333333433333333333333;
		rom_data[110] <= 3840'h7777777665555554544434433333333233357ACCCECECECCCB9988AA99998888788A9999998898654432489A98888888888777754202234567766665577778877766676666665555886666555544346BCCA8532232323232332323233333333333323332333333333323333233233233333233333323333333333334788875434343000000000000000000000000000000234333434343433433433343333433433434343444344444344434434343443433334333333333333333333434334343433334344455555555555555555656667677666555443322222222022222022222222233333333343334333333888888887777777665555554544434433333333233357ACCCECECECCCB9988AA99998888788A9999998898654432489A98888888888777754202234567766665577778877766676666665555886666555544346BCCA8532232323232332323233333333333323332333333333323333233233233333233333323333333333334788875434343000000000000000000000000000000234333434343433433433343333433433434343444344444344434434343443433334333333333333333333434334343433334344455555555555555555656667677666555443322222222022222022222222233333333343334333333;
		rom_data[111] <= 3840'h77777776655555554444433333333323322347ACCCCECCBAAA999AAAA98887888899998999999865542358A9988888888887765542222345666677776777777777777666676555579855655554543347CEEEB854323223233233333323323332333333333333333333333233323323332333333333333333333333677555533434332200000000000000000000000000023333334343334333433343333433343443444344444443444444443444434343343333433333333343343433434343443433343444545555555555555556666667766655544332222220222202022202020222333333434334334343338888887777777776655555554444433333333323322347ACCCCECCBAAA999AAAA98887888899998999999865542358A9988888888887765542222345666677776777777777777666676555579855655554543347CEEEB85432322323323333332332333233333333333333333333323332332333233333333333333333333367755553343433220000000000000000000000000002333333434333433343334333343334344344434444444344444444344443434334333343333333334334343343434344343334344454555555555555555666666776665554433222222022220202220202022233333343433433434333;
		rom_data[112] <= 3840'h7777766666555554544434433333333323323479BCCCBA88899ABBAA998877788888888889999875533468888877787667767755543345567666777767777665566567667776665887566555554443347ACEEEC975332232323323333333333333333333333233323332333233333333323333333333333323335785445444433333222000000000000000000000000233433434334343434434343343433434343443444444444444444444444434434343434333334334333333434343443444433334344455555555555555556666667767655543332222202202022220202020202223334334333433433343888887777777766666555554544434433333333323323479BCCCBA88899ABBAA998877788888888889999875533468888877787667767755543345567666777767777665566567667776665887566555554443347ACEEEC975332232323323333333333333333333333233323332333233333333323333333333333323335785445444433333222000000000000000000000000233433434334343434434343343433434343443444444444444444444444434434343434333334334333333434343443444433334344455555555555555556666667767655543332222202202022220202020202223334334333433433343;
		rom_data[113] <= 3840'h77777666555555544444433333333332332323468ACCB9889ABBBBA9998767788987777889899986543477888876676556667755555567766656777777776666665677767888876776777555555443435579BCEECA8653322323332332333233333333333333332333233233323233233333333333333332345557543444444434332200000000000000000000000003443433434434343433434343434343434344344444444444444444444444443434343343434333333343433434344444344343343444444555555555555566667766766555433322202202220200020200002022233334433443433343338888878777777666555555544444433333333332332323468ACCB9889ABBBBA9998767788987777889899986543477888876676556667755555567766656777777776666665677767888876776777555555443435579BCEECA865332232333233233323333333333333333233323323332323323333333333333333234555754344444443433220000000000000000000000000344343343443434343343434343434343434434444444444444444444444444343434334343433333334343343434444434434334344444455555555555556666776676655543332220220222020002020000202223333443344343334333;
		rom_data[114] <= 3840'h777766665555554544443443333333333323223458BCBA889BCCCA9888875678888775678888888755457778887667666566765555566775556777888877666767777776788888877777765555554444444579BCEECBA87543232323333333333333333333333333333333323333233333333333333332335896554344544444333322000000000000000000000002334343434343444343443434343434434344444444444444444444444444444444434334343343434343333434344434444344343343444555555555555556676777766655543332222200200202020000000020222233334443433434343488878777777766665555554544443443333333333323223458BCBA889BCCCA9888875678888775678888888755457778887667666566765555566775556777888877666767777776788888877777765555554444444579BCEECBA875432323233333333333333333333333333333333233332333333333333333323358965543445444443333220000000000000000000000023343434343434443434434343434344343444444444444444444444444444444444343343433434343433334343444344443443433434445555555555555566767777666555433322222002002020200000000202222333344434334343434;
		rom_data[115] <= 3840'h7777666555555545444434333333332323323323368AAAA9ACCCB98887755777788766577777888776778777887666765555665566566766678888888777667777777677889899877877765555555444433445689ACEECCA98653323232333323333333323333333233233333323333323333333333323478A744433454343333332220000000000000000000000034434343433444344434343443444343443434434444444454444444444444443434343434343434333343434344434444444434333444454454444554555566676777765554433222000200200000000000000022223333444343443434343888877777777666555555545444434333333332323323323368AAAA9ACCCB98887755777788766577777888776778777887666765555665566566766678888888777667777777677889899877877765555555444433445689ACEECCA98653323232333323333333323333333233233333323333323333333333323478A744433454343333332220000000000000000000000034434343433444344434343443444343443434434444444454444444444444443434343434343434333343434344434444444434333444454454444554555566676777765554433222000200200000000000000022223333444343443434343;
		rom_data[116] <= 3840'h777766655555554444434343333333333232323233568888ACCB98887555557778876667877788887888887777775555556666666666777778988888777677777787656888998887776566556555555544443334568ACCCCECBA8555333232333333333333333333333332333333333333333333323356898653343443433333222202000000000000000000000244433443434343443434444434443444434444444444444544445444444444444444444434343434343434343434344444344444434333444544444445455555667777776555443322222000000000000000000002022233343444434434343488887777777766655555554444434343333333333232323233568888ACCB98887555557778876667877788887888887777775555556666666666777778988888777677777787656888998887776566556555555544443334568ACCCCECBA85553332323333333333333333333333323333333333333333333233568986533434434333332222020000000000000000000002444334434343434434344444344434444344444444444445444454444444444444444444343434343434343434343444443444444343334445444444454555556677777765554433222220000000000000000000020222333434444344343434;
		rom_data[117] <= 3840'h7776665555555454444434333333332323332332323345568AB9877754434567788877788888888778899877888766655677776777767778889988877777777777755568899888765555555556676665545443333445789BCCECCCBA8654333332333323333333333333333323332333332333333456899754333434333333222000020000000000000000000023443434444444444344434344444444434434444444444454454544454544444444343434443443443434343434444444444444444434344445444444444555566777767666554433220000000000000000000000202223333444344443444444887777777776665555555454444434333333332323332332323345568AB9877754434567788877788888888778899877888766655677776777767778889988877777777777755568899888765555555556676665545443333445789BCCECCCBA8654333332333323333333333333333323332333332333333456899754333434333333222000020000000000000000000023443434444444444344434344444444434434444444444454454544454544444444343434443443443434343434444444444444444434344445444444444555566777767666554433220000000000000000000000202223333444344443444444;
		rom_data[118] <= 3840'h77766665555555444443433333333333323233233323333468987776433345777888788888888877679BB988898888767887666677677678888888877677887788755678888877765434556667666554445554444443456789ABCCEEECB97554433323333333333333333333333332333333333467889875444334333333332020200000000000000000000002454443443443434444434444434444344434444444444454454545455544544444444444443443443444343434434444444444444444434344444343344444555567777776655544322220200000000000000000000222223333444443444434348877777777766665555555444443433333333333323233233323333468987776433345777888788888888877679BB988898888767887666677677678888888877677887788755678888877765434556667666554445554444443456789ABCCEEECB9755443332333333333333333333333333233333333346788987544433433333333202020000000000000000000000245444344344343444443444443444434443444444444445445454545554454444444444444344344344434343443444444444444444443434444434334444455556777777665554432222020000000000000000000022222333344444344443434;
		rom_data[119] <= 3840'h77666655555554444434343333333333333233332333233345775665434457888888778888888876789ABA99999988888987755776666678888888777778877877666778887766554345577655444333333344445544434456778ABCCCECBA988654333333333333333333233333333333433458BA866554544333333332222000000000000000000000000033444344434444444444444444444444444444444444544454545454554455445444444444344434444434443443444444444444444444434343443433443445555667777776655443332020000000000000000000000202223334444444444344447877777777666655555554444434343333333333333233332333233345775665434457888888778888888876789ABA99999988888987755776666678888888777778877877666778887766554345577655444333333344445544434456778ABCCCECBA988654333333333333333333233333333333433458BA86655454433333333222200000000000000000000000003344434443444444444444444444444444444444444454445454545455445544544444444434443444443444344344444444444444444443434344343344344555566777777665544333202000000000000000000000020222333444444444434444;
		rom_data[120] <= 3840'h7776665555554544444434343333332332332323333233323444555567567899888776789898877888888889AA999889AA98755666776787777777766677788877777778887655444455655433333323232323345555555545555778ABBCCCCCCBA877543323333333333333333333335775568B9655444344432322223020000000000000000000000000234344443444344444444444444444444444444444444544554555545545545455454544444444444434444344434444444444444444444444343434333333444555666777776655544432220200000000000000000000000222333344444444444444877777777776665555554544444434343333332332332323333233323444555567567899888776789898877888888889AA999889AA98755666776787777777766677788877777778887655444455655433333323232323345555555545555778ABBCCCCCCBA877543323333333333333333333335775568B9655444344432322223020000000000000000000000000234344443444344444444444444444444444444444444544554555545545545455454544444444444434444344434444444444444444444444343434333333444555666777776655544432220200000000000000000000000222333344444444444444;
		rom_data[121] <= 3840'h6766656555555444444343333333333332323333232332333233334589888899888877789AA98888876556789999989ABBA987567776678876555555555677775557787767765565555543323232323232323232333456555565555556899ABCCCCCCBA8654433233333323332333235787557875444444433222202222000000000000000000000000002333443444444444444444444444444444444444444445455545555455555455554544544444444444444444444444444444454444445454443433333333334344455566777766555544332222000000000000000000000002222333444444444444444777777776766656555555444444343333333333332323333232332333233334589888899888877789AA98888876556789999989ABBA987567776678876555555555677775557787767765565555543323232323232323232333456555565555556899ABCCCCCCBA8654433233333323332333235787557875444444433222202222000000000000000000000000002333443444444444444444444444444444444444444445455545555455555455554544544444444444444444444444444444454444445454443433333333334344455566777766555544332222000000000000000000000002222333444444444444444;
		rom_data[122] <= 3840'h7766655555555444444343433333333333332323333323333332333479878899989888889999877765555555789989ABBBA998777755778775434455556567654445566566655555443333232333233323332323323344444577675544557789AABBBBBBA98875533332333333333478754555554444333333222222020000000000000000000000000223444434434444444444444444444444444444444445454554555555555555555455455454544444444444444444344444444444454454454444344333333333444455566677665554443332222020000000000000000000000222233344444444444444787777777766655555555444444343433333333333332323333323333332333479878899989888889999877765555555789989ABBBA998777755778775434455556567654445566566655555443333232333233323332323323344444577675544557789AABBBBBBA98875533332333333333478754555554444333333222222020000000000000000000000000223444434434444444444444444444444444444444445454554555555555555555455455454544444444444444444344444444444454454454444344333333333444455566677665554443332222020000000000000000000000222233344444444444444;
		rom_data[123] <= 3840'h7666655555554444444434333333332332323333232333232332332356656788999898999887555445677554578999AAAA98987675556777654344555555665555456665555444433333233323323323323233232332333334456776555455566778899AABCCCA9775543332333336BA534554443333323232222200200000000000000000002300000344444344444444444444444545454545454444545454554555555555555555555555554545444444444444444444444444444454544454544443433333333333344455566666555544433332222020000000000000000000002022333444444445445444777777777666655555554444444434333333332332323333232333232332332356656788999898999887555445677554578999AAAA98987675556777654344555555665555456665555444433333233323323323323233232332333334456776555455566778899AABCCCA9775543332333336BA534554443333323232222200200000000000000000002300000344444344444444444444444545454545454444545454554555555555555555555555554545444444444444444444444444444454544454544443433333333333344455566666555544433332222020000000000000000000002022333444444445445444;
		rom_data[124] <= 3840'h66656555555545444434334333333332333323233333233332333333334445567788989987543333456777545689A9A9A988776677655555544444444555555555555555433333333332332333332332332332333233232333344555555555555555567789ABCCCCBB987553332358A84344433333322222222000200000000000000000000000002234444344444444444445454544544454544545454545454554555555555555555555555555454544454544444444444444444544454454545454434333332323333344555655555554433333232222020000000000000000000002222333444454545454547777777766656555555545444434334333333332333323233333233332333333334445567788989987543333456777545689A9A9A988776677655555544444444555555555555555433333333332332333332332332332333233232333344555555555555555567789ABCCCCBB987553332358A8434443333332222222200020000000000000000000000000223444434444444444444545454454445454454545454545455455555555555555555555555545454445454444444444444444454445445454545443433333232333334455565555555443333323222202000000000000000000000222233344445454545454;
		rom_data[125] <= 3840'h66665555555444444444343333333333323233332323333323332333333334445556777775322333455567755578AAA999876556776544445444443434333334554444333333323233233233323333333233233233323333333333334445454555544455567789AACCCCB987654489633334332323220200000000000000000000000000000000033443434444444444444454454445454554545454554545555555555555555555555555555554554545444544544444445444454545445454545544443333333333333345555555555443333222222220200200000000000000000022223333444445454545457777777766665555555444444444343333333333323233332323333323332333333334445556777775322333455567755578AAA999876556776544445444443434333334554444333333323233233233323333333233233233323333333333334445454555544455567789AACCCCB98765448963333433232322020000000000000000000000000000000003344343444444444444445445444545455454545455454555555555555555555555555555555455454544454454444444544445454544545454554444333333333333334555555555544333322222222020020000000000000000002222333344444545454545;
		rom_data[126] <= 3840'h666665555555544444443434333333333333332333323323333333232333332333344444433223343444467644578AA98875555555544333333333333332332323323232333333333333333333333233333233233233333333333333333434445665544444545557889AABBAA978873202233322222020202000000000000000000000000000003444443444444444444444445455454554545555455545445555555555555555555555555555555545454545454454545444454545545454545545553433323232323334445555555444433322222220202020000000000000000002022222333444545454545477777767666665555555544444443434333333333333332333323323333333232333332333344444433223343444467644578AA98875555555544333333333333332332323323232333333333333333333333233333233233233333333333333333434445665544444545557889AABBAA9788732022333222220202020000000000000000000000000000034444434444444444444444454554545545455554555454455555555555555555555555555555555454545454544545454444545455454545455455534333232323233344455555554444333222222202020200000000000000000020222223334445454545454;
		rom_data[127] <= 3840'h666565555545544444343434333333323232323323233333332333333332333323332333333233333333456532358887755434333333333333333333232333333333333333333323333323333333333323333233233333333333333333333334555455665544444445557889BBB9842000222222220222000000000000000000000000000000023434344444444444445454545554555545555455555555555455555555555555555555555555554554545454544544544454545445455554555455544333322322232334455555554443333222222222202020200000000000000002022222333444455455455477777776666565555545544444343434333333323232323323233333332333333332333323332333333233333333456532358887755434333333333333333333232333333333333333333323333323333333333323333233233333333333333333333334555455665544444445557889BBB98420002222222202220000000000000000000000000000000234343444444444444454545455545555455554555555555554555555555555555555555555555545545454545445445444545454454555545554555443333223222323344555555544433332222222222020202000000000000000020222223334444554554554;
		rom_data[128] <= 3840'h6665555555554444444444334333333333333323333333323333333333333333333333323233233332333444333456554333333333333333333333333333333333233333333333333333333332333333333333233332333333333333343434433443456777555544433445568A997300222222222202020200000000000000000000000000000344434344444444444544544555555545555555555555555555555555555555555555555555555555555545545545455445445454555555555555555443333322222233344555554544333323222222202222202202000000000002002022222334444455455545777777676665555555554444444444334333333333333323333333323333333333333333333333323233233332333444333456554333333333333333333333333333333333233333333333333333333332333333333333233332333333333333343434433443456777555544433445568A997300222222222202020200000000000000000000000000000344434344444444444544544555555545555555555555555555555555555555555555555555555555555545545545455445445454555555555555555443333322222233344555554544333323222222202222202202000000000002002022222334444455455545;
		rom_data[129] <= 3840'h6656555555554544444434343333333332332333233333333333333333333333333333333333332333333333333334333333333333333333333323333333323333333333333333333333333333333333333333332333333333343434333434334434344555555665544333347AAA7300202220020002000020000000000000000000000000002434444444444454545455455555555555555555555555555555555555555555555555555555555555555455455455454454545455554555555555555443332222222233344455554444333222222222222222222022022020000020020222222333444545555555777776766656555555554544444434343333333332332333233333333333333333333333333333333333332333333333333334333333333333333333333323333333323333333333333333333333333333333333333333332333333333343434333434334434344555555665544333347AAA7300202220020002000020000000000000000000000000002434444444444454545455455555555555555555555555555555555555555555555555555555555555555455455455454454545455554555555555555443332222222233344455554444333222222222222222222022022020000020020222222333444545555555;
		rom_data[130] <= 3840'h6655555555555444444443433433333333333323333332333333333333333333333333333333233333233333333333333333332333333333333333333333333333333333333333333333333333333333333333333333333333333333443434343343434344445566555553338CEB7322220222200000000232000000000000000000000000024443344444445454544545545554555555555555555555555555555555555555555555555555555555555555545555544555455455455555555555555443323222222223344455454443333232222222222222222222222202222002002002222333444455555545777776666655555555555444444443433433333333333323333332333333333333333333333333333333233333233333333333333333332333333333333333333333333333333333333333333333333333333333333333333333333333333333443434343343434344445566555553338CEB7322220222200000000232000000000000000000000000024443344444445454544545545554555555555555555555555555555555555555555555555555555555555555545555544555455455455555555555555443323222222223344455454443333232222222222222222222222202222002002002222333444455555545;
		rom_data[131] <= 3840'h6665555555555545444443434333333333333333323333333333333333333333333333333333332333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333334334343434343434343434343344444556776558CC84323202200200000000354200000000000000000000000245444444444444454545555555555555555555555555555555555555555555555555555555555555555555555555455545454545545555555555555555443332222222233334454544443333232323223333323323222222222202220220222222333344545555555777767666665555555555545444443434333333333333333323333333333333333333333333333333333332333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333334334343434343434343434343344444556776558CC84323202200200000000354200000000000000000000000245444444444444454545555555555555555555555555555555555555555555555555555555555555555555555555455545454545545555555555555555443332222222233334454544443333232323223333323323222222222202220220222222333344545555555;
		rom_data[132] <= 3840'h656555555555455454444444334333333233323333333333333333333333333333333333332333333333333333333333333333333333333333333333333323333333333333333333333333333333333333333333333333333343343433434343444344444343434344557755575322222220000000000003872000000000000000000000003544444444444454454545545555555555555555555555555555555555555555555555555555555555555555555555555554554554554555555555555554433322222022233444444444443333323323333333333333333232322222222220222222333444555555557777766665655555555545545444444433433333323332333333333333333333333333333333333333233333333333333333333333333333333333333333333333332333333333333333333333333333333333333333333333333333334334343343434344434444434343434455775557532222222000000000000387200000000000000000000000354444444444445445454554555555555555555555555555555555555555555555555555555555555555555555555555555455455455455555555555555443332222202223344444444444333332332333333333333333323232222222222022222233344455555555;
		rom_data[133] <= 3840'h666555555555554544444434343333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333433343333333333333333333333333434344343443443443434444344343445554322000220200000000000002662000000000000000000000025544444444444454554555555555555555555555555555555555555555555555555555555555555555555555555555555455555545555555555555555554433222202222233344444444433333333333333334334333333333332322222222222223233444555555557777666666655555555555454444443434333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333343334333333333333333333333333343434434344344344343444434434344555432200022020000000000000266200000000000000000000002554444444444445455455555555555555555555555555555555555555555555555555555555555555555555555555555545555554555555555555555555443322220222223334444444443333333333333333433433333333333232222222222222323344455555555;
		rom_data[134] <= 3840'h665655555555455545444444434343333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333343333343343333433333333333333333334343434343434444344444344443443443444334333220200002000000000000000220000000000000000000000245534444444444545555555555555555555555555555555555555555555555555555555555555555555555555555555555554555555555555555555555554443322222022233334444444444343343434344444444444444343333333332222222222333344455555557776766666565555555545554544444443434333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333334333334334333343333333333333333333434343434343444434444434444344344344433433322020000200000000000000022000000000000000000000024553444444444454555555555555555555555555555555555555555555555555555555555555555555555555555555555555455555555555555555555555444332222202223333444444444434334343434444444444444434333333333222222222233334445555555;
		rom_data[135] <= 3840'h665555555555554454444443343433333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333343333434333433443334343333434333333334343343434434344434344444344444444444443432332220020000000000000000000000000000000000000002575444444444555455555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555443332220222233343444444444444444444454555455545444444443333333323222223233444555555557677766666555555555555445444444334343333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333334333343433343344333434333343433333333434334343443434443434444434444444444444343233222002000000000000000000000000000000000000000257544444444455545555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555544333222022223334344444444444444444445455545554544444444333333332322222323344455555555;
		rom_data[136] <= 3840'h656555555555555544544444434333333333333333333333333333333333333333333333333333333333333333333333333333333433333333434333333333333333343334343333343343343433334343343333333433333434343444443444443444444444444443444433452220000000000000000000000000000000000000000003785444445454445555555555555555555555555555555555555555555555555555555655555555555555555555555555555555555555555555555555555555443333222202223343444445444444454444555555555555555545444444433333323222333344555555557777666665655555555555554454444443433333333333333333333333333333333333333333333333333333333333333333333333333333343333333343433333333333333334333434333334334334343333434334333333343333343434344444344444344444444444444344443345222000000000000000000000000000000000000000000378544444545444555555555555555555555555555555555555555555555555555555565555555555555555555555555555555555555555555555555555555544333322220222334344444544444445444455555555555555554544444443333332322233334455555555;
		rom_data[137] <= 3840'h665655555555555455444444443433333333333333333333333333333333434333343333333333333333333333433333334343433334343434333343333333343433334333433443433434343434434343433433433344343443444434444444444444444444444444444433542200000000000000000000000000000000000000000036764444445455555555555555555555555555555555555555555555555555555555565655556555555555555555555555555555555555555555555555555555544333322222223333444454454545555555555555555555555555555545444433333333333444555555557767666666565555555555545544444444343333333333333333333333333333333343433334333333333333333333333343333333434343333434343433334333333334343333433343344343343434343443434343343343334434344344443444444444444444444444444444443354220000000000000000000000000000000000000000003676444444545555555555555555555555555555555555555555555555555555555556565555655555555555555555555555555555555555555555555555555554433332222222333344445445454555555555555555555555555555554544443333333333344455555555;
		rom_data[138] <= 3840'h666665555555555555454444444443433333333333333333333343333333333434333433333333333333333343334343433333334333333343343433434333333334343434334333443334343434343434343434334333444344443444444444444444444444444444444433320000000000000000000000000000000000000000002355554444454554545555555555555555555555555555555555555555555555555555565565665665655555555555555555555555555555555555555555555555544433332222223333444454545455555555555656566665555555555555555544443333333444555555557776766666666555555555555545444444444343333333333333333333334333333333343433343333333333333333334333434343333333433333334334343343433333333434343433433344333434343434343434343433433344434444344444444444444444444444444444443332000000000000000000000000000000000000000000235555444445455454555555555555555555555555555555555555555555555555555556556566566565555555555555555555555555555555555555555555555554443333222222333344445454545555555555565656666555555555555555554444333333344455555555;
		rom_data[139] <= 3840'h665655555555555554544544443434333333333333333333333333433434334333433333433333333333434343433433343343433434344434433343333343344343333434343444344443434434434444343433434344434443444444444444444444444444444444444432220000000000000000000000000000000000000000024555444444545545555555555555555555555555555555555555555555555555555565566565655656555555555555555555555555555555555555555555555555554433332222223334344454545455555555556566666666666666656656565555544433334445555555557777666666565555555555555454454444343433333333333333333333333343343433433343333343333333333343434343343334334343343434443443334333334334434333343434344434444343443443444434343343434443444344444444444444444444444444444444443222000000000000000000000000000000000000000002455544444454554555555555555555555555555555555555555555555555555555556556656565565655555555555555555555555555555555555555555555555555443333222222333434445454545555555555656666666666666665665656555554443333444555555555;
		rom_data[140] <= 3840'h666665555555555555454444444343434333333333333333333433343333433344334343334343334343334343443434334343434334334343434343443334334343443433434343443434443443444434434344343443444344444444444444444444444445454444444442000000000000000000000000233222000000000000245544444545455555555555555555555555555555555555555555556565565565666656566666665566565556555555555555555555555555555555555555555555555444333232232333444455555555555555656666666666766667777777776665555544444445555555557777666666666555555555555545444444434343433333333333333333343334333343334433434333434333434333434344343433434343433433434343434344333433434344343343434344343444344344443443434434344344434444444444444444444444444545444444444200000000000000000000000023322200000000000024554444454545555555555555555555555555555555555555555555656556556566665656666666556656555655555555555555555555555555555555555555555555544433323223233344445555555555555565666666666676666777777777666555554444444555555555;
		rom_data[141] <= 3840'h665656555555555554554544444434333433333333343434343334333434343433434333433334343434443434434434343434334343434343434343433434343434434344344344434444344444434344444434343444444444444444444444444444444544544545444442200000000000000000000003577532000000000002235544545454555555555555555555555555555565555565656565656656565656565666665666656566565655655555555555555555555555555555555555565655555544333332323333444555545555555555566666666677677777777777777777665555444454555555557776666666565655555555555455454444443433343333333334343434333433343434343343433343333434343444343443443434343433434343434343434343343434343443434434434443444434444443434444443434344444444444444444444444444444454454454544444220000000000000000000000357753200000000000223554454545455555555555555555555555555556555556565656565665656565656566666566665656656565565555555555555555555555555555555555556565555554433333232333344455554555555555556666666667767777777777777777766555544445455555555;
		rom_data[142] <= 3840'h666565655555555555554544444443443343433434333333334343343343434344344343343434334343434443443434443434343443434344434434343434434344344443444443444344443434344443443444344434344444444444444444445454545454545444444444322000000000000000000034579754000000000002245545454545555555555555555555555555555556556566565656556666666665666566566666666666665566565555555555555555555555555555555555566565655554443333333333444555555555555556566666666667677777777777888887776555555545555555557777776666656565555555555555454444444344334343343433333333434334334343434434434334343433434343444344343444343434344343434443443434343443434434444344444344434444343434444344344434443434444444444444444444545454545454544444444432200000000000000000003457975400000000000224554545454555555555555555555555555555555655656656565655666666666566656656666666666666556656555555555555555555555555555555555556656565555444333333333344455555555555555656666666666767777777777788888777655555554555555555;
		rom_data[143] <= 3840'h666665655555555555554554444444434334343434344344343343434334334343433443434334343444444344434443434434344343443443434343434344344444443444434444444444444444444444434444444344444444444444444454454454544545454445454555543220000000000000000245568875200000000000355554545555555555555555555555555555556665656566666666666666666666656665666666666656556665655655555555555555555555555555555555656666665555443333333334445555555555555555666666666676777777778788888888887765555455555555557777676666666565555555555555455444444443433434343434434434334343433433434343344343433434344444434443444343443434434344344343434343434434444444344443444444444444444444444443444444434444444444444444445445445454454545444545455554322000000000000000024556887520000000000035555454555555555555555555555555555555666565656666666666666666666665666566666666665655666565565555555555555555555555555555555565666666555544333333333444555555555555555566666666667677777777878888888888776555545555555555;
		rom_data[144] <= 3840'h666666555555555555455455544444434343434334343434334343433434344344344344434443443434444444444444443444443444344443444344434443443434444444444444444444444444444444444444434444444444444444444544545454445455455454544555433202000000000000000355458A850000000000035865545555555555555555555555555656556565656565656566666666666666666666666666666666666666665655555555655555555555555555565565656566566665555444333333344445555555555555556566656666677777777888888889888887765555555555655577777677666666555555555555455455544444434343434334343434334343433434344344344344434443443434444444444444443444443444344443444344434443443434444444444444444444444444444444444444434444444444444444444544545454445455455454544555433202000000000000000355458A8500000000000358655455555555555555555555555556565565656565656565666666666666666666666666666666666666666656555555556555555555555555555655656565665666655554443333333444455555555555555565666566666777777778888888898888877655555555556555;
		rom_data[145] <= 3840'h666666656555555555555554444444343434343434344434343444344343434443443443444434344444444444444444344434434434444444434443444444444444444444444444444444444444444444444444444444444445444545455445445545545554545545454543322200000000000000004454546873000200000025886545555555555555555555555555555656565666666566666666666666666666666666666666666666666656656656555555555555555555555555655666666666666555544443333334445555555555555555555656665666777777788888899999988887765555555656567777676766666665655555555555555444444434343434343434443434344434434343444344344344443434444444444444444434443443443444444443444344444444444444444444444444444444444444444444444444444444444544454545544544554554555454554545454332220000000000000000445454687300020000002588654555555555555555555555555555565656566666656666666666666666666666666666666666666666665665665655555555555555555555555565566666666666655554444333333444555555555555555555565666566677777778888889999998888776555555565656;
		rom_data[146] <= 3840'h666666665555555555555555454444443434343443434344444343443444344344444344434344443444444444444444444444444444444444444444444444444444444444444444444444544544444444444444444444444544545445444554555455455455555455545542200200000000000000035555555553022222220257765555555555555555555555555565666565656666656666666666666666666666766666666666666666666666666665666655656565656555565666566656656666667655554444434344445555555555555555565565556666667777888889999999998888766555555665657777777766666666555555555555555545444444343434344343434444434344344434434444434443434444344444444444444444444444444444444444444444444444444444444444444444444454454444444444444444444444454454544544455455545545545555545554554220020000000000000003555555555302222222025776555555555555555555555555556566656565666665666666666666666666666676666666666666666666666666666566665565656565655556566656665665666666765555444443434444555555555555555556556555666666777788888999999999888876655555566565;
		rom_data[147] <= 3840'h6666666655555555555554554544444344343434343434434344444344344344343444434444434444444444444444444444444444444444444444444444444444444444444444454454454444454444454444444444444444544545454554554545545545545555554555430200000000000000000355554455532233323346776555555555555555555555555666566566666666666666666666666666666666666666666666666666667666666666666565656555555556555565666656666666666667655544443344444555555555555555556555555565666777777888889999AAAA998877666555556656777767676666666655555555555554554544444344343434343434434344444344344344343444434444434444444444444444444444444444444444444444444444444444444444444444454454454444454444454444444444444444544545454554554545545545545555554555430200000000000000000355554455532233323346776555555555555555555555555666566566666666666666666666666666666666666666666666666666667666666666666565656555555556555565666656666666666667655544443344444555555555555555556555555565666777777888889999AAAA998877666555556656;
		rom_data[148] <= 3840'h766666566565555555555555545444443444344344344344443434344443443444444444344344344444444444444444444444444444444444444444444444444444444544444444454544454544454545444444444444545455454554554554555555555555545555545553200000000000000000035555555685432322345775555555555555555555555555556565665656566666666656666666666666666766666666766667666666666666666665666666566665665555556566666666666666666766555544444444555555555555555565555555555565666777788889999AAAAAA9988777655556666677776777766666566565555555555555545444443444344344344344443434344443443444444444344344344444444444444444444444444444444444444444444444444444444544444444454544454544454545444444444444545455454554554554555555555555545555545553200000000000000000035555555685432322345775555555555555555555555555556565665656566666666656666666666666666766666666766667666666666666666665666666566665665555556566666666666666666766555544444444555555555555555565555555555565666777788889999AAAAAA99887776555566666;
		rom_data[149] <= 3840'h66666666565555555555555545444444444344344344444344444444344444443444444444444444444444454545454544444444444444444444444444444444444444444554545454545454545545454545545454444444554555545554555555555555555555555555555422000000000000000024555555578753322245565555555555555555555555556656666666666666666666666666677676767676766777666666666676676666676676666666665666565656666665656666666666666666667655554444444545555555555555555565555555555566677777888889AAABBBAA99887777655566657777776766666666565555555555555545444444444344344344444344444444344444443444444444444444444444454545454544444444444444444444444444444444444444444554545454545454545545454545545454444444554555545554555555555555555555555555555422000000000000000024555555578753322245565555555555555555555555556656666666666666666666666666677676767676766777666666666676676666676676666666665666565656666665656666666666666666667655554444444545555555555555555565555555555566677777888889AAABBBAA9988777765556665;
		rom_data[150] <= 3840'h777666666556555555555555455454444344434444434444444444444444434444434444444444444444454445444544545454545445454444444444444444454544445455454545454545545545455455554544454545454555455554555554555555555555555555555554222000000000000000355555555687532224555555555555555555555555656566665666666666666666666666667667676767676777767776666676677767667676766666666666566656665565656666666666666667777767655554545455555555555555555565555555555555667676777888899AABBBBBA99887776656666677777776777666666556555555555555455454444344434444434444444444444444434444434444444444444444454445444544545454545445454444444444444444454544445455454545454545545545455455554544454545454555455554555554555555555555555555555554222000000000000000355555555687532224555555555555555555555555656566665666666666666666666666667667676767676777767776666676677767667676766666666666566656665565656666666666666667777767655554545455555555555555555565555555555555667676777888899AABBBBBA998877766566666;
		rom_data[151] <= 3840'h767666665655555555555555554544444443444434444344444444444443444444444444444444444445454554545454454545454454544545454444444444445445455545554555545555555555545555455454544545555554555555555555555555555555555555555554220000000000000000455555555578643357765555555555555555555556566665666666666666666666666667776776777677777767767676777667776666777676766666666666666565566666666666666666666676766677665555555555555555555555555555555555555556556666667788899AABBBCBBA9988777666666677777777767666665655555555555555554544444443444434444344444444444443444444444444444444444445454554545454454545454454544545454444444444445445455545554555545555555555545555455454544545555554555555555555555555555555555555555554220000000000000000455555555578643357765555555555555555555556566665666666666666666666666667776776777677777767767676777667776666777676766666666666666565566666666666666666666676766677665555555555555555555555555555555555555556556666667788899AABBBCBBA99887776666666;
		rom_data[152] <= 3840'h766666666565655555555555555554444444344444444444444444444444444444444444444444544444545454555455455555455545454545454545454545454545454555455555555555555555555555555555555455455555555555555555555555555555555555555554222000000000000024555555555558876776655555555555555555555556666666666666666677766777776667667767776767777777776777767776767777767777676666666666666666666566666666666666666666767767766555555555555555555555555555555555555555555655566778899AABBBBBBBA988777766666677777777766666666565655555555555555554444444344444444444444444444444444444444444444444544444545454555455455555455545454545454545454545454545454555455555555555555555555555555555555455455555555555555555555555555555555555555554222000000000000024555555555558876776655555555555555555555556666666666666666677766777776667667767776767777777776777767776767777767777676666666666666666666566666666666666666666767767766555555555555555555555555555555555555555555655566778899AABBBBBBBA9887777666666;
		rom_data[153] <= 3840'h776766666566556555555555555445444444444444444444444444444444444444444444444444445454545545555554554555555455454544545445445454454554555555555555555555555555555555555554555555555555555555555555555555555555555555555554320020000000000355555555555557888875555555555555555555555556666666666666676666666766677777677777777777777777777777777777777777777677676767676666666666666666666666666766676777777677766655555555555555555555555555555555555555555555556777899AABBBBBBBA988877776666777777776776766666566556555555555555445444444444444444444444444444444444444444444444444445454545545555554554555555455454544545445445454454554555555555555555555555555555555555554555555555555555555555555555555555555555555555554320020000000000355555555555557888875555555555555555555555556666666666666676666666766677777677777777777777777777777777777777777777677676767676666666666666666666666666766676777777677766655555555555555555555555555555555555555555555556777899AABBBBBBBA9888777766667;
		rom_data[154] <= 3840'h676666666655665555555555555554544444444444444444444444444444444444444444545454544545455455545555555555555555554545454554554545455455455555555555555555555555555555555555545555455555555545555555555555555555555555555554322000000000003455555555555555677655555555555555555556665555666666555555656667777767766777767777777777777777777777777777777777777777776767676766666666666666666666676676767777777777776655555555555555555555555555555555555555555555555677899AABBBBBBBA998887776766677777777676666666655665555555555555554544444444444444444444444444444444444444444545454544545455455545555555555555555554545454554554545455455455555555555555555555555555555555555545555455555555545555555555555555555555555555554322000000000003455555555555555677655555555555555555556665555666666555555656667777767766777767777777777777777777777777777777777777777776767676766666666666666666666676676767777777777776655555555555555555555555555555555555555555555555677899AABBBBBBBA9988877767666;
		rom_data[155] <= 3840'h776676666656656555555555555554545444444444444444444444545444444454544454454544545455554555555555555555555555555555555545545455555555555555555555555555555555555555555454434344333444345676544555555555555555555555555554320220000000034555555555555555555555555555555565444679ACCB755555689ABBBAA97655677776777777777777777777777777777777777777777777777777777776776676766666676666676766767677777777777777777665555555555555555555555555555555555555555555555668889AABABAAAAA998888777667777777777776676666656656555555555555554545444444444444444444444545444444454544454454544545455554555555555555555555555555555555545545455555555555555555555555555555555555555555454434344333444345676544555555555555555555555555554320220000000034555555555555555555555555555555565444679ACCB755555689ABBBAA97655677776777777777777777777777777777777777777777777777777777776776676766666676666676766767677777777777777777665555555555555555555555555555555555555555555555668889AABABAAAAA9988887776677;
		rom_data[156] <= 3840'h7776666666665565555555555555554545444444444444445454545445444454544545454554554545455555555555555555555555555555555555554555554555555555555555555555555555555545555545558ABA758CBBB989BBBBBA7544555555555555555555555554222022000002355555555555555555555555655555556554589AA988BEEA76889AABCCCCEEEEC86567777777777777777777777777777777777777777777777777777777777676777676666666666666676767677777777777777776555555555555555454555555555555555555555554455556778899AAAAAAA999988887777666776777767776666666665565555555555555554545444444444444445454545445444454544545454554554545455555555555555555555555555555555555554555554555555555555555555555555555555545555545558ABA758CBBB989BBBBBA7544555555555555555555555554222022000002355555555555555555555555655555556554589AA988BEEA76889AABCCCCEEEEC86567777777777777777777777777777777777777777777777777777777777676777676666666666666676767677777777777777776555555555555555454555555555555555555555554455556778899AAAAAAA999988887777666;
		rom_data[157] <= 3840'h6666766666666655555555555555555454444444444444544445445444545445445454554545454555555555555555555555555555555555555555555555555555555555555555555555555555555665545689AACEECCCCEEEECBCCCBCCECA76766555555555555555555554220200000003555555555555555555565556556565655558BB9997558EEB88BB9877788889BEEEC9767777777777777777777777777777777777777777777777777777777777777777767777777776776767767777777777777777766555555555555444545445455555555555555544444555557788899AAAAA9989888877777677767767776666766666666655555555555555555454444444444444544445445444545445445454554545454555555555555555555555555555555555555555555555555555555555555555555555555555555665545689AACEECCCCEEEECBCCCBCCECA76766555555555555555555554220200000003555555555555555555565556556565655558BB9997558EEB88BB9877788889BEEEC9767777777777777777777777777777777777777777777777777777777777777777767777777776776767767777777777777777766555555555555444545445455555555555555544444555557788899AAAAA9989888877777677;
		rom_data[158] <= 3840'h7676766666666665655555555555555554554454545454445545454454454545455555455455454545455555555555555555555555555555555555555555555555555555555555555555555556788ACA878BCEEECCCEEEEECECCCECCCCCCEECBBCAAA999998889A88777787754322200002555555555555555555566656666665566558AC98877569ECB99CEBA9888878777BEECA866766777777777777777777777777777777777777777777777777777777677777776777677777776777777777777777777776665555555545444444445454545555455545444444444555677788899A9A99888877777777777777777677676766666666665655555555555555554554454545454445545454454454545455555455455454545455555555555555555555555555555555555555555555555555555555555555555555556788ACA878BCEEECCCEEEEECECCCECCCCCCEECBBCAAA999998889A88777787754322200002555555555555555555566656666665566558AC98877569ECB99CEBA9888878777BEECA866766777777777777777777777777777777777777777777777777777777677777776777677777776777777777777777777776665555555545444444445454545555455545444444444555677788899A9A99888877777777777;
		rom_data[159] <= 3840'h6766767666666665555555555555555555544554545454554554545545455454554555555555554555555555555555555555555555555555555555555555555555555555555555555555555579BCCEEECCCEEECCECECEEECECCEECEEEEEEEEEEEEEEEEEEEEEEEEEEECCCCCBBA986533223345555555555555556565555555655666568AAA9BCBAAACCCCCACEEEBBCECCCB98ACCCCA8899877777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777665555544444444444444454544444444444444444444455557778889999998888777777777777777776776766767666666665555555555555555555544554545454554554545545455454554555555555554555555555555555555555555555555555555555555555555555555555555555555555555579BCCEEECCCEEECCECECEEECECCEECEEEEEEEEEEEEEEEEEEEEEEEEEEECCCCCBBA986533223345555555555555556565555555655666568AAA9BCBAAACCCCCACEEEBBCECCCB98ACCCCA8899877777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777665555544444444444444454544444444444444444444455557778889999998888777777777777;
		rom_data[160] <= 3840'h76767766666666656555555555555555545554545545554554554554554545554555555555555555555555555555555555555555555555555555555555555555555555555555555555555667CCECCCCEEEECCCCCECCCCCECECECECECEECECEEEEEEEEEEEEEEEEEEEEEEEEEECECECB9877975677776667775556555545555555565578889ABEEEEECCBABCCCEECACCEEEEEEEEEECECCCEEB767777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777776655554444444444444444444444444444444434434444555567788889998888777667677777777777676776767766666666656555555555555555545554545545554554554554554545554555555555555555555555555555555555555555555555555555555555555555555555555555555555555667CCECCCCEEEECCCCCECCCCCECECECECECEECECEEEEEEEEEEEEEEEEEEEEEEEEEECECECB9877975677776667775556555545555555565578889ABEEEEECCBABCCCEECACCEEEEEEEEEECECCCEEB76777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777665555444444444444444444444444444444443443444455556778888999888877766767777777;
		rom_data[161] <= 3840'h7777666666666666665555555555555555555555545545554555554554555545554555555555555555555555555555555555555555555555555555555555555555555555555555555568ACCEEEECCCEECCCCCCBCCCCCCCCCCCCCCCCCCCCCCEEEEECEECCCEEEEEEEEEEEEEEEEEECCCBC99CE858AAAAA77AB97764455355676556656787679889BEEECC97899EEEEEEEEEEEEEEEEEEEEEEEC86677777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777655555443343433434444444443433333333333333434445557788888899987777666666677777777777767777666666666666665555555555555555555555545545554555554554555545554555555555555555555555555555555555555555555555555555555555555555555555555555555568ACCEEEECCCEECCCCCCBCCCCCCCCCCCCCCCCCCCCCCEEEEECEECCCEEEEEEEEEEEEEEEEEECCCBC99CE858AAAAA77AB97764455355676556656787679889BEEECC97899EEEEEEEEEEEEEEEEEEEEEEEC86677777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777655555443343433434444444443433333333333333434445557788888899987777666666677777;
		rom_data[162] <= 3840'h677676766666666565665555555555555555545455455545555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555556899ACCECECCECEEEECECCCCCBABAABBCCCBCBCCCBBBCCCCCECBCECECCEEECEEEECEEEEEEEEEEEEECBECA9987788AAAA98ABAA8789898778988788667778A9668A8CABB86778ABBA9BCC878BEEEEEEEEEEEEEA8778999887787777777778777777777777777777777777777777777777777777777777777777777777777777777666555444433433334344444433333333333323333333445556778888898988877766566667777777777667677676766666666565665555555555555555545455455545555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555556899ACCECECCECEEEECECCCCCBABAABBCCCBCBCCCBBBCCCCCECBCECECCEEECEEEECEEEEEEEEEEEEECBECA9987788AAAA98ABAA8789898778988788667778A9668A8CABB86778ABBA9BCC878BEEEEEEEEEEEEEA87789998877877777777787777777777777777777777777777777777777777777777777777777777777777777776665554444334333343444444333333333333233333334455567788888989888777665666677777;
		rom_data[163] <= 3840'h7677667676666656665555555555555555555555555555555555555555555555555555555555555555555555555555555565555555555555555555555555555555688888889BCCCCCEEEEEEEEEEEEEEEECCBBCCCCBBBCECCCBCCCBBBBCCBCA89CBBBBBBB998ACB9A99CEEBCEEEEEEBCCCCCEEEEEEEECECECBBBCCCECBABBA9999888899988988979BCCA75569A8898AEE84458AEEEECEEEEEEEEAABCECBCCBBBB98777777777777777777777777777777777777777777777777777777777777777777777777777665544433333333334343443333333333323232333344455666788899998887776665666677777777777767677667676666656665555555555555555555555555555555555555555555555555555555555555555555555555555555565555555555555555555555555555555688888889BCCCCCEEEEEEEEEEEEEEEECCBBCCCCBBBCECCCBCCCBBBBCCBCA89CBBBBBBB998ACB9A99CEEBCEEEEEEBCCCCCEEEEEEEECECECBBBCCCECBABBA9999888899988988979BCCA75569A8898AEE84458AEEEECEEEEEEEEAABCECBCCBBBB98777777777777777777777777777777777777777777777777777777777777777777777777777665544433333333334343443333333333323232333344455666788899998887776665666677777;
		rom_data[164] <= 3840'h7776776766666666666565555555555555555555555555555555555555555555555555555555555555555555555555556555656555656656555555555577655558CECBCCCBCCEEEEEEEEEEEEEEEEEEEEEECCEEEEECCCCCECBECBBBBBCBCCBA9899BAA7677565777757CEECAABCBBBABCCCCEEEEEEEEEEECEEEEEEEEEECCCCCBABBCCCCCAACB88A98899CC98579877789EC97535EEEEEEEEEEEEEEEEECECEEEEEEEECA8777777777777777777777777777777777777777777777777777777777777777777777776655544433332333333434434333333323222222233344455666778899988888766665566677777777777777776776766666666666565555555555555555555555555555555555555555555555555555555555555555555555555556555656555656656555555555577655558CECBCCCBCCEEEEEEEEEEEEEEEEEEEEEECCEEEEECCCCCECBECBBBBBCBCCBA9899BAA7677565777757CEECAABCBBBABCCCCEEEEEEEEEEECEEEEEEEEEECCCCCBABBCCCCCAACB88A98899CC98579877789EC97535EEEEEEEEEEEEEEEEECECEEEEEEEECA8777777777777777777777777777777777777777777777777777777777777777777777776655544433332333333434434333333323222222233344455666778899988888766665566677777;
		rom_data[165] <= 3840'h7777667677666666665656555555555555555555555555555555555555555555555555555555555555555555555556565656556565656565655555458BBBAA88ACCECCECCCEEEEEEEEEEEEEEEEEEEEEEEEEEEEECCCCCBCBBAB99ABBBCBBCCCBAA9AAA97544555555568CEEC9679A9BECEECEAACEEEEEEECCCEEEEEEEEEECCBABBBCEECEECACC88876789BEE887887889CCCBBABEEEEEEEEEEEEEEEEEEEECB88CEEEEEE877787777777777777777777777777777777777777777777777777777777777777777777655544333223223333343333333333232222232333344555667777889998888776555666777777777777777777667677666666665656555555555555555555555555555555555555555555555555555555555555555555555556565656556565656565655555458BBBAA88ACCECCECCCEEEEEEEEEEEEEEEEEEEEEEEEEEEEECCCCCBCBBAB99ABBBCBBCCCBAA9AAA97544555555568CEEC9679A9BECEECEAACEEEEEEECCCEEEEEEEEEECCBABBBCEECEECACC88876789BEE887887889CCCBBABEEEEEEEEEEEEEEEEEEEECB88CEEEEEE877787777777777777777777777777777777777777777777777777777777777777777777655544333223223333343333333333232222232333344555667777889998888776555666777777;
		rom_data[166] <= 3840'h767777676766666666665555555555555555555555555555555555555555555555555555555555555555555555555555565656566656656566555569CCCCECECCECCCCCCEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEBBBCCCBBBBBCBAABCBCCBCBBBABBCB9A977887755554578ACCCBECAECB999978ACCEECCEECBAACCCCCCCBABACCCCECCCEEEAACC77875688AC9655789A9BBCCCABEEEC9888889CEEEEEEEEECC98BEEEEEEA777777777777777777777777777777777777777777777777777777777777777777777665544333222222223333333333332332222222323334455566677788888988877555566777777777777676767777676766666666665555555555555555555555555555555555555555555555555555555555555555555555555555565656566656656566555569CCCCECECCECCCCCCEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEBBBCCCBBBBBCBAABCBCCBCBBBABBCB9A977887755554578ACCCBECAECB999978ACCEECCEECBAACCCCCCCBABACCCCECCCEEEAACC77875688AC9655789A9BBCCCABEEEC9888889CEEEEEEEEECC98BEEEEEEA7777777777777777777777777777777777777777777777777777777777777777777776655443332222222233333333333323322222223233344555666777888889888775555667777777;
		rom_data[167] <= 3840'h7777777776766666666566665555555555555555555555555555555555555555555555555555555555555555655566666566666666666666655677AECCCCECECCECCCCCEEEEEEEEEEEEEEEEEEEEECCEEEEEEEECBABCBBBCCCCCCABAABBCCAAABBCCCAABBCECBA9987765557ACCCA8887777778888888ABA9867CBBAABB889BCCEEECCEEBCC9BEB889757779A754578889AA9A99CEEE977655557BEEEEEEEEEEBABACEEEEB777787777777777777777777777777777777777777777777777777777777777777776555443322222222323333333333333222232333333445555566777888898888876555666777777777777777777777776766666666566665555555555555555555555555555555555555555555555555555555555555555655566666566666666666666655677AECCCCECECCECCCCCEEEEEEEEEEEEEEEEEEEEECCEEEEEEEECBABCBBBCCCCCCABAABBCCAAABBCCCAABBCECBA9987765557ACCCA8887777778888888ABA9867CBBAABB889BCCEEECCEEBCC9BEB889757779A754578889AA9A99CEEE977655557BEEEEEEEEEEBABACEEEEB777787777777777777777777777777777777777777777777777777777777777777776555443322222222323333333333333222232333333445555566777888898888876555666777777;
		rom_data[168] <= 3840'h77777777776776666665656566655555555555555555555555555555555555555555555555555555555555656556565666666666666666655689CCEEECCECCCCECCCECEEEEEEEEEEEEEEEEEECCCCCCCEEEEEEEECCCCCCCECCCBBBA99BBCBBCCCCBBBBCCCCEECECEEECA85556777764358977788887788877757BABBBA98789BBEEEEEECBECC99CB799877789A97667788899ACCCEEEECCA89776778CEEEEEEEEEB8BCCEEEA777787777777777777777777777777777777777777777777777777777777777777765554333222022222323333333323332323233333444455555666677888888888765555677777787777777777777777776776666665656566655555555555555555555555555555555555555555555555555555555555656556565666666666666666655689CCEEECCECCCCECCCECEEEEEEEEEEEEEEEEEECCCCCCCEEEEEEEECCCCCCCECCCBBBA99BBCBBCCCCBBBBCCCCEECECEEECA85556777764358977788887788877757BABBBA98789BBEEEEEECBECC99CB799877789A97667788899ACCCEEEECCA89776778CEEEEEEEEEB8BCCEEEA77778777777777777777777777777777777777777777777777777777777777777776555433322202222232333333332333232323333344445555566667788888888876555567777778;
		rom_data[169] <= 3840'h777777776777676666666666656555555555555555555555555555555555555555555555555555555555555665656666566666666666655558BEEECEECECCCECCCCEEEEEEEEEEEEEEEEEECBAAAAABCCCCEEEEEEECECEEECCCCABBBAAABCBBCCCBBABBBBCCCBBBBCCECCA889AA989865579A9888ABBBB98899769BBBCAAA8888A9BCCCEECCCA888C988898878AA97778778ABA9ACEECEEEE9CCCC9657BCEECCEEEEBCCCBEEE8877777777777777777777777777777777777777777777777777777777777777766555443323222202222223232323333333333333334445555556667778888988887665666777788877777777777777776777676666666666656555555555555555555555555555555555555555555555555555555555555665656666566666666666655558BEEECEECECCCECCCCEEEEEEEEEEEEEEEEEECBAAAAABCCCCEEEEEEECECEEECCCCABBBAAABCBBCCCBBABBBBCCCBBBBCCECCA889AA989865579A9888ABBBB98899769BBBCAAA8888A9BCCCEECCCA888C988898878AA97778778ABA9ACEECEEEE9CCCC9657BCEECCEEEEBCCCBEEE88777777777777777777777777777777777777777777777777777777777777777665554433232222022222232323233333333333333344455555566677788889888876656667777888;
		rom_data[170] <= 3840'h77777777776767666666656566665655555555555555555555555555555555555555555555555555556556565665665666666666665665578CEEEEEECCCCEECCCCCCEEEEEEEECEECEEECCBAABAABBCCCCCECCEEEEEECCCCBB9ABBBBBABECABCBABBBAACCCCBBBA9ABCCCCCCEECCCEEC7579A898889BCA999AA89BAABBAA99888755778A88877778878AAA88777899855567ABB9AAECAEE84689EEE96977EECEEEEEEECBBCECB9877777777777777777777777777777777777777777777777777777777777776555544333222020202222232323333333333333333345555555666677788888887765666677788887777777777777777776767666666656566665655555555555555555555555555555555555555555555555555556556565665665666666666665665578CEEEEEECCCCEECCCCCCEEEEEEEECEECEEECCBAABAABBCCCCCECCEEEEEECCCCBB9ABBBBBABECABCBABBBAACCCCBBBA9ABCCCCCCEECCCEEC7579A898889BCA999AA89BAABBAA99888755778A88877778878AAA88777899855567ABB9AAECAEE84689EEE96977EECEEEEEEECBBCECB987777777777777777777777777777777777777777777777777777777777777655554433322202020222223232333333333333333334555555566667778888888776566667778888;
		rom_data[171] <= 3840'h777777777776766766666666666566565655555555555555555555555555555555555555555565555555555566666666666666665568ACEEEEEEECCCBCEEEBBCEECCCCCCEEECECCECCCCCA9ABAABAAACCBCCCEEEECCCCCBAAABAABCBBBC99BBCCBCBCBCCCCCCBCCB9CCCA889AEECEBAC96AB9ACEECCBBCCABA99AACC98978989B9A9757755567888876788775558BA6655678989A8CCBCB778889CEEE857CEEEEEEEEEECABBCCB877777777777777777777777777777777777777777777777777777777777765554433322202020220222223233333433444443444455555555666677788888877666677778888877777777777777777776766766666666666566565655555555555555555555555555555555555555555565555555555566666666666666665568ACEEEEEEECCCBCEEEBBCEECCCCCCEEECECCECCCCCA9ABAABAAACCBCCCEEEECCCCCBAAABAABCBBBC99BBCCBCBCBCCCCCCBCCB9CCCA889AEECEBAC96AB9ACEECCBBCCABA99AACC98978989B9A9757755567888876788775558BA6655678989A8CCBCB778889CEEE857CEEEEEEEEEECABBCCB8777777777777777777777777777777777777777777777777777777777777655544333222020202202222232333334334444434444555555556666777888888776666777788888;
		rom_data[172] <= 3840'h777777777777777776666666666666666556565555556565555555555555555555555555555556555656666666666666666666568AEEEEEEEEECECCCCCECBCCEEECCCBEEEECCCCCB9ABCA9AAABBBBBBCBACCCCCECCCEECBBAAA999BBAAA9AABBBBBBCCBBBBBAAEEECABAA98999ABA999A98AA88A99CCCCBBAA8889C99AA999BCECCB999A9888888A988887777767888567777779887BCCEE998898CECEC9BEEEEEEEEEEEEECCECBA9777777777777777777777777777777777777777777777777777777777655544333222200000002022222223333333444444344455555555566677778887777665677778888877777777777777777777777776666666666666666556565555556565555555555555555555555555555556555656666666666666666666568AEEEEEEEEECECCCCCECBCCEEECCCBEEEECCCCCB9ABCA9AAABBBBBBCBACCCCCECCCEECBBAAA999BBAAA9AABBBBBBCCBBBBBAAEEECABAA98999ABA999A98AA88A99CCCCBBAA8889C99AA999BCECCB999A9888888A988887777767888567777779887BCCEE998898CECEC9BEEEEEEEEEEEEECCECBA97777777777777777777777777777777777777777777777777777777776555443332222000000020222222233333334444443444555555555666777788877776656777788888;
		rom_data[173] <= 3840'h7777777777776766766666666666656556565656555555565555555556555555555656555555555565566565656666666676568CECBBCEEEEECCCBBCBCBBCCECECCCCEEEECBBCBABA9ABBBBBCBBBAAAAACCCCCECBCCCCBBBAAAAAABA99AAAAAABBBBBABCCBCABBBBBAA988887678889BBBA9BA9BAABCBB9899A89BCBBB9888ACECB99ABCBAAAAA99A9888876776778A867876778887ACCEEC988778A89AABCEEEEEEEEEEEEEEEEEEECB98777777777777777777777777777777777777777777777777777665554433332220002020202022223333334344444444445555555555566667777777766666777778888777777777777777777776766766666666666656556565656555555565555555556555555555656555555555565566565656666666676568CECBBCEEEEECCCBBCBCBBCCECECCCCEEEECBBCBABA9ABBBBBCBBBAAAAACCCCCECBCCCCBBBAAAAAABA99AAAAAABBBBBABCCBCABBBBBAA988887678889BBBA9BA9BAABCBB9899A89BCBBB9888ACECB99ABCBAAAAA99A9888876776778A867876778887ACCEEC988778A89AABCEEEEEEEEEEEEEEEEEEECB98777777777777777777777777777777777777777777777777777665554433332220002020202022223333334344444444445555555555566667777777766666777778888;
		rom_data[174] <= 3840'h77777777777777776767666666666666666565565656566565655556656565655565556556556555556566666666666667557ACCAABEEEEEECCBBBBBBBABEEEEEEEEEEEECAACCBABBBBBBBCBCBBAAABCCEECEECCBBBBAABAACCCCBBAAAB9ABBBBAAABBCCCCCCCA88AAB9888766876678BB99ABABBBCAA988BC889CECBBBA989988999AAABAABBA9ABA888887778878BC78878989ABAABACEECA888878ABAAACEEEEEEEEEECEEEEEEEECECA976677777777777777777777777777777777777777777777766555443332222020000000000202222333334334444444455555555555666777777766555566778778887777777777777777777777776767666666666666666565565656566565655556656565655565556556556555556566666666666667557ACCAABEEEEEECCBBBBBBBABEEEEEEEEEEEECAACCBABBBBBBBCBCBBAAABCCEECEECCBBBBAABAACCCCBBAAAB9ABBBBAAABBCCCCCCCA88AAB9888766876678BB99ABABBBCAA988BC889CECBBBA989988999AAABAABBA9ABA888887778878BC78878989ABAABACEECA888878ABAAACEEEEEEEEEECEEEEEEEECECA97667777777777777777777777777777777777777777777776655544333222202000000000020222233333433444444445555555555566677777776655556677877888;
		rom_data[175] <= 3840'h7777777777777777777666766666666666666665666666565565666565665555555565556566565566566566666666766558CEB89CEEEEEECCBBCCCBBAAEEEEEEEEEEECAAABBBABCEBBBBBCCCCCAABCEECCEEECBABBBABBAACEECCBABAABBBBB9AAABBCCBCCCB9889CCCBBA98999777789A9CBBCCCCA8A98AA8ABCCCA9BCB9998AB9998AAAACCAABAAA9A998756568888989CB89ACC988ACCEEA8ABCCABCBAACEEEEEEECCBCEEEEEEEEEEEECA76777777777777777777777777777777777777777777776555443333222000000000000002222232333334444454554545555555556677776656555555677778788777777777777777777777777777666766666666666666665666666565565666565665555555565556566565566566566666666766558CEB89CEEEEEECCBBCCCBBAAEEEEEEEEEEECAAABBBABCEBBBBBCCCCCAABCEECCEEECBABBBABBAACEECCBABAABBBBB9AAABBCCBCCCB9889CCCBBA98999777789A9CBBCCCCA8A98AA8ABCCCA9BCB9998AB9998AAAACCAABAAA9A998756568888989CB89ACC988ACCEEA8ABCCABCBAACEEEEEEECCBCEEEEEEEEEEEECA76777777777777777777777777777777777777777777776555443333222000000000000002222232333334444454554545555555556677776656555555677778788;
		rom_data[176] <= 3840'h777777777777776776777776666666666665666666666666666665666666655656565565555656655565666666676765679EEA8AEEEEEEECBBCCCCBBAABEEEEEEEEEB9AABAABABACBAABABBABBCBCCECCCCCCCCABCCBBBAAABECBAABAABCCBB99ABAABCBAAEBAA98BBCCEECAABAA998889A9ABCCBBA99C98888ACCCCB88CCBACCCB88899889CCABB99A9888A965457867999BA9A89CA779A8ACEBACEC9ACCB9ACCBEEEECECA8AEEEEEEEEEEEEC877777777777777777777777777777777777777877776555444333222202000000000000002222333333334444544545455555555667777655555555567777787877777777777777777777776776777776666666666665666666666666666665666666655656565565555656655565666666676765679EEA8AEEEEEEECBBCCCCBBAABEEEEEEEEEB9AABAABABACBAABABBABBCBCCECCCCCCCCABCCBBBAAABECBAABAABCCBB99ABAABCBAAEBAA98BBCCEECAABAA998889A9ABCCBBA99C98888ACCCCB88CCBACCCB88899889CCABB99A9888A965457867999BA9A89CA779A8ACEBACEC9ACCB9ACCBEEEECECA8AEEEEEEEEEEEEC8777777777777777777777777777777777777778777765554443332222020000000000000022223333333344445445454555555556677776555555555677777878;
		rom_data[177] <= 3840'h7777777777777777777767666666666666666666666665666665665656656665665656566665565666666666667676679CEEC9CEEEEEEECCCCCCBBBAABCEEEEEECCB99ABA9AABBA99ABAABAAABBBCCBCCCBCCCBABCCBABAAAABB99AAAABBBB999CCA9BCC9ACBAA88BBABEEEAABA9AA9A99B9889AABBAAC988888ABCCEAABCCCBBA889999889BC999A998778ACB8668C9578888A978CCA879889CEBAA9ABBBBA9AA99CEEEEEC87BB89EEEEEEEEEEB87777777777777777777777777777777788888777765554433322202000000000000020220222333333434444454444555555566677776655555555667777777777777777777777777777777777767666666666666666666666665666665665656656665665656566665565666666666667676679CEEC9CEEEEEEECCCCCCBBBAABCEEEEEECCB99ABA9AABBA99ABAABAAABBBCCBCCCBCCCBABCCBABAAAABB99AAAABBBB999CCA9BCC9ACBAA88BBABEEEAABA9AA9A99B9889AABBAAC988888ABCCEAABCCCBBA889999889BC999A998778ACB8668C9578888A978CCA879889CEBAA9ABBBBA9AA99CEEEEEC87BB89EEEEEEEEEEB87777777777777777777777777777777788888777765554433322202000000000000020220222333333434444454444555555566677776655555555667777777;
		rom_data[178] <= 3840'h77777777777777777677767666666776666666666666666666666666666666665665666665665565656566666666568CEEECEEEEEEEEEECCCBBBBAAAACEEECCCBBBA9AAABBCBABCA99BBBBBBBBBCCCBBBCCCCBBBCCBAA9AAAAAAA999AAAAA999BBB8ACECCC9A988ACCABCCCABEEBABAA88A98888CEEEAB9878989CECEEECCCE99A9899998ABBA888ABB9888ACEECBCEC768A98778BACE977797ACECCC9AABBBBBBA99CEEEEEC9A98AEEEECBBCEEEC87777777777777777777777777777777888887777555443332222002000000000000000222222233433334444444454555555666667665555555555677777777777777777777777777777777677767666666776666666666666666666666666666666665665666665665565656566666666568CEEECEEEEEEEEEECCCBBBBAAAACEEECCCBBBA9AAABBCBABCA99BBBBBBBBBCCCBBBCCCCBBBCCBAA9AAAAAAA999AAAAA999BBB8ACECCC9A988ACCABCCCABEEBABAA88A98888CEEEAB9878989CECEEECCCE99A9899998ABBA888ABB9888ACEECBCEC768A98778BACE977797ACECCC9AABBBBBBA99CEEEEEC9A98AEEEECBBCEEEC8777777777777777777777777777777788888777755544333222200200000000000000022222223343333444444445455555566666766555555555567777777;
		rom_data[179] <= 3840'h7777777777777777777776767676676676666767666666666666666666665666665665565665666666666666666669EEEEEEEEEEEEEECCCCAABBAAAABCCCCCABCAA9AABBCCCBAAAA9ABCCCBCCBBCCBBCCCBBABBBCCBAA9AAAAAABA99AAB999A9AB99ACCABCCA999BCECEECBCCECCBA9888A989999CEE99A88778BCBCECBCCCB98888889A99AAA8888ABBA999ABCCCCB998A887679B99CB7666777878CB99BBBBABBBA9CCCCEECBABEEBECCECBCEEEC877777777777777777777777777778888888777665544332222000000000000000002020222232333333344444455555555566666665555445555567777777777777777777777777777777777776767676676676666767666666666666666666665666665665565665666666666666666669EEEEEEEEEEEEEECCCCAABBAAAABCCCCCABCAA9AABBCCCBAAAA9ABCCCBCCBBCCBBCCCBBABBBCCBAA9AAAAAABA99AAB999A9AB99ACCABCCA999BCECEECBCCECCBA9888A989999CEE99A88778BCBCECBCCCB98888889A99AAA8888ABBA999ABCCCCB998A887679B99CB7666777878CB99BBBBABBBA9CCCCEECBABEEBECCECBCEEEC877777777777777777777777777778888888777665544332222000000000000000002020222232333333344444455555555566666665555445555567777777;
		rom_data[180] <= 3840'h77777777777777777777776767677676767666767666666666666666656666565666666666666666666666666656BEEEEEEEEEEEEECCECCBBBBAABBCCECBBAAABAA99AABCCA9999AABBBBBCCBAACCCCCCCBAABBBCCA999ABBBBAAAAAAA999AA999999BA9AAECA8ABACCCBBABEECA89A98889A99878A99AB877799BBACECCCCA988779999867887CB888ABA9656788666468867877A9ABB87677689AAACB99BBBBBBBAABCCBABBBBCEECCAAEECEEEEEB877777777777777777777777777888888887766554433222202000000000000000002022222232333333344545555455555566666555544445555677777777777777777777777777777777777776767677676767666767666666666666666656666565666666666666666666666666656BEEEEEEEEEEEEECCECCBBBBAABBCCECBBAAABAA99AABCCA9999AABBBBBCCBAACCCCCCCBAABBBCCA999ABBBBAAAAAAA999AA999999BA9AAECA8ABACCCBBABEECA89A98889A99878A99AB877799BBACECCCCA988779999867887CB888ABA9656788666468867877A9ABB87677689AAACB99BBBBBBBAABCCBABBBBCEECCAAEECEEEEEB87777777777777777777777777788888888776655443322220200000000000000000202222223233333334454555545555556666655554444555567777777;
		rom_data[181] <= 3840'h7777777777777777777776776777667677666767667666666666666666666666666565656666566656566666656BEEEEEEEEEEEEEECEBBBCBAAAACCCCCCC9ABBCBAABBBBBAAAAA999AAAABBABCEECBBBCCCAABBBAA999AAAA99999AAA9ABBAA99899889BBA889A98677755679CCCBC88889999978BB888A9755558A9CCBBA9876558887857ACB9BE99AA889854345556887668888BCBB98888ACCB87CCCB9AAAABAABBABCCBBCBABCEEECCEEEEEEEEC87777777777777777777777777888888888776655543322200000000000000000000020202222222333344445555555555565666555554444555567777777777777777777777777777777777776776777667677666767667666666666666666666666666565656666566656566666656BEEEEEEEEEEEEEECEBBBCBAAAACCCCCCC9ABBCBAABBBBBAAAAA999AAAABBABCEECBBBCCCAABBBAA999AAAA99999AAA9ABBAA99899889BBA889A98677755679CCCBC88889999978BB888A9755558A9CCBBA9876558887857ACB9BE99AA889854345556887668888BCBB98888ACCB87CCCB9AAAABAABBABCCBBCBABCEEECCEEEEEEEEC87777777777777777777777777888888888776655543322200000000000000000000020202222222333344445555555555565666555554444555567777777;
		rom_data[182] <= 3840'h777777777777777777777777776776677676767677677666666666666666666666666666656666666666666666AEEEEEEEEEEEEEECCCCBBCBBABCCCCBABBABCBAAAAABCBABBBB99AA99A9AAABCCCCBBCCCCCCBBB9AA99AAA999999AAAA999AA99989888999899AA87777788899CCCCA8888879CBBCC8779976433578998765555789887769CCCA9BC9888999754457789877678788998658899BEC8789CBAAAAABABAAAAACBCCEECBCEEEEEEECEEEC98877777777777777777777777888888888877655544322222000000000000000000002022222222223334445555555555555555555555444455556677777777777777777777777777777777777777776776677676767677677666666666666666666666666666656666666666666666AEEEEEEEEEEEEEECCCCBBCBBABCCCCBABBABCBAAAAABCBABBBB99AA99A9AAABCCCCBBCCCCCCBBB9AA99AAA999999AAAA999AA99989888999899AA87777788899CCCCA8888879CBBCC8779976433578998765555789887769CCCA9BC9888999754457789877678788998658899BEC8789CBAAAAABABAAAAACBCCEECBCEEEEEEECEEEC988777777777777777777777778888888888776555443222220000000000000000000020222222222233344455555555555555555555554444555566777777;
		rom_data[183] <= 3840'h777777777777777777777777777767777777776767676766666666666666666666666666666666666666666668EEEEEEEEEEEEECCCCBCBCBBAABCBBBB9AABBA999ABABCBBCBCB9AA99AABCBBBBCBAABCCBCECBBC9ABAAAAAA9999AAAAA9BBB98988988889989AA99899BBAAA99CCBB9889887ACEAACA7799985445465554455668BA98778BB9CCB8BA8799999788888887787577877766667888ACB877B99CBAABBBABBA9BBAABEECCCCEEEEEEACCC98777777777777777777777778888888888777655543332200000000000000000000002020222222223334445555555555555555555554444455566677777777777777777777777777777777777777777767777777776767676766666666666666666666666666666666666666666668EEEEEEEEEEEEECCCCBCBCBBAABCBBBB9AABBA999ABABCBBCBCB9AA99AABCBBBBCBAABCCBCECBBC9ABAAAAAA9999AAAAA9BBB98988988889989AA99899BBAAA99CCBB9889887ACEAACA7799985445465554455668BA98778BB9CCB8BA8799999788888887787577877766667888ACB877B99CBAABBBABBA9BBAABEECCCCEEEEEEACCC987777777777777777777777788888888887776555433322000000000000000000000020202222222233344455555555555555555555544444555666777777;
		rom_data[184] <= 3840'h77777777777777777777777777777777777767776767676777776666666666666666666666666666666666656AEEEEEEEEEEEEECECBBBBBBBAABCBBBA99AAAA989A9AABCCBAAA9AAABCCEECCCCBAAABBBABCCBBBABCB99AA9A9AABBAA9CCCBA888899988999AAABA99ABC99A9ABB88788988899B98BB88AAB9766667555557777ACA87999A88CCC87878888988A98778777A9657787778A876788ACA79CA8998ABBAABBA9AA9999BCCCCCCCCEECCEEC976777777777777777777777888888888877655543332220200000000000000000000002220222222233345555555555555555555555555455556677777777777777777777777777777777777777777777777777767776767676777776666666666666666666666666666666666656AEEEEEEEEEEEEECECBBBBBBBAABCBBBA99AAAA989A9AABCCBAAA9AAABCCEECCCCBAAABBBABCCBBBABCB99AA9A9AABBAA9CCCBA888899988999AAABA99ABC99A9ABB88788988899B98BB88AAB9766667555557777ACA87999A88CCC87878888988A98778777A9657787778A876788ACA79CA8998ABBAABBA9AA9999BCCCCCCCCEECCEEC97677777777777777777777788888888887765554333222020000000000000000000000222022222223334555555555555555555555555545555667777777;
		rom_data[185] <= 3840'h77777777777777777777777777777777777777777777776767676667666666666666666666666656666667657BEEEEEEEEEEEEECCCCCCAABBBBBBBA9999A9A99989AA9ABBA9A9ABCCECEECEEECCBAABBAAACCBB9BBBB98888ABBBBAA89BCCBAA8889998899ABBAAA8999BB989AA878999887878AA89C9889A8788777788888878AB867999988BC975678888989A98777788AA87767889AA9755789A97BBC9779ABB9AABAA9AAA988ACECCECEEEEEEEEC86677777777777777777777888888888777655443322220000000000000000000000202022222222233444555565555554455555555555555566777787887777777777777777777777777777777777777777777777777777776767676667666666666666666666666656666667657BEEEEEEEEEEEEECCCCCCAABBBBBBBA9999A9A99989AA9ABBA9A9ABCCECEECEEECCBAABBAAACCBB9BBBB98888ABBBBAA89BCCBAA8889998899ABBAAA8999BB989AA878999887878AA89C9889A8788777788888878AB867999988BC975678888989A98777788AA87767889AA9755789A97BBC9779ABB9AABAA9AAA988ACECCECEEEEEEEEC8667777777777777777777788888888877765544332222000000000000000000000020202222222223344455556555555445555555555555556677778788;
		rom_data[186] <= 3840'h77777777777777777777777777777777777777777777767677767666666666666666666666666666666666668CEEEEEEEEEECACECCCCCAABBBBBBA9A999A988989ABA9999AABCCCEEEECCEEEECBBBABAABCCCBAABBABA8789ABCBABA889AA8AC989988899BABA9988BBACC989A889BCB987667AAA98A86689888865578AA8888887578989AABCA5458AA999AABC98998889A99A87789B978975788887B8BEA9B9ABAABBAAABB99999ACCECEEEEEECECEC9777777777777777777778888888877776554433322020000000000000000000000020220222222233344555566555554444555555555555667778788887777777777777777777777777777777777777777777777777777767677767666666666666666666666666666666666668CEEEEEEEEEECACECCCCCAABBBBBBA9A999A988989ABA9999AABCCCEEEECCEEEECBBBABAABCCCBAABBABA8789ABCBABA889AA8AC989988899BABA9988BBACC989A889BCB987667AAA98A86689888865578AA8888887578989AABCA5458AA999AABC98998889A99A87789B978975788887B8BEA9B9ABAABBAAABB99999ACCECEEEEEECECEC977777777777777777777888888887777655443332202000000000000000000000002022022222223334455556655555444455555555555566777878888;
		rom_data[187] <= 3840'h7777777777777777777777777777777777777777777777676777767777766666666666666666656666666568CEEEEEEEEEEEE8BCCBAAAABBBBBBB99BB99A999ABB99A99889A9BCECECECECECCCAABCC9BBBBBBAAABABCBAAB9AAAABB989998898999999998AAABA9BCC98BA999989BCCBA8857BB9997558BB87886678888779B97778989BBBA87579AAA988BCCA8898888AB99BA988AC978AA766787599ACEB989AAABBAAAAA99AAA9ABCEECEEEBEECEEEE9877777777777777777878888787777555433322220000000000000000000000000202222222232334455566555554444445555555555667777778888777777777777777777777777777777777777777777777777777777676777767777766666666666666666656666666568CEEEEEEEEEEEE8BCCBAAAABBBBBBB99BB99A999ABB99A99889A9BCECECECECECCCAABCC9BBBBBBAAABABCBAAB9AAAABB989998898999999998AAABA9BCC98BA999989BCCBA8857BB9997558BB87886678888779B97778989BBBA87579AAA988BCCA8898888AB99BA988AC978AA766787599ACEB989AAABBAAAAA99AAA9ABCEECEEEBEECEEEE9877777777777777777878888787777555433322220000000000000000000000000202222222232334455566555554444445555555555667777778888;
		rom_data[188] <= 3840'h777777777777777777777777777777777777777777777777767677777776666666666666565666566666669EEEEEEEEEEEEEE9CCBBBA9ABBBCBAA99A99999BA9A989A9989A99CCCBCECCECEECBAABAABBBAAA9AAA988899AAAAAACCAA888AA978ABA9A9988BCEC9888A999889889BEEE9898679AAA8658A8875566777789889AC9778778988756788999997AEEBAA998878988AA9778887799888AA76788AAAAAA99AABA9AA9AA9AAA9ABBECCCBABEEEEECCB8777777777777777878888877776555433322202000000000000000000000000002002022222333445556655554544444455555555566777788888877777777777777777777777777777777777777777777777777777777767677777776666666666666565666566666669EEEEEEEEEEEEEE9CCBBBA9ABBBCBAA99A99999BA9A989A9989A99CCCBCECCECEECBAABAABBBAAA9AAA988899AAAAAACCAA888AA978ABA9A9988BCEC9888A999889889BEEE9898679AAA8658A8875566777789889AC9778778988756788999997AEEBAA998878988AA9778887799888AA76788AAAAAA99AABA9AA9AA9AAA9ABBECCCBABEEEEECCB87777777777777778788888777765554333222020000000000000000000000000020020222223334455566555545444444555555555667777888888;
		rom_data[189] <= 3840'h77777777777777777777777777777777777777777777777777777676767666666666666566666656666668EEEEEEEEEEEEEEECECBBAAABBBBBBBABA99A99BCAA9889A999AA9ABCCBCCCCECCCCBAA9AAABBAAA9ABBA888AABB99A9AAA9878778789CAA9AA9BCECCBA989898888857BEECA8887779AA856BB9888777777888777887788777875566888889977ACCBBAABC87888899A778888776798AB77755668AACCECB99999ABAABA99BABCECCCCEECEECBCEB76677777777777777887877776555443322220200000000000000000000000000202022222223344556555554444344445455555566677788888887777777777777777777777777777777777777777777777777777777777777676767666666666666566666656666668EEEEEEEEEEEEEEECECBBAAABBBBBBBABA99A99BCAA9889A999AA9ABCCBCCCCECCCCBAA9AAABBAAA9ABBA888AABB99A9AAA9878778789CAA9AA9BCECCBA989898888857BEECA8887779AA856BB9888777777888777887788777875566888889977ACCBBAABC87888899A778888776798AB77755668AACCECB99999ABAABA99BABCECCCCEECEECBCEB7667777777777777788787777655544332222020000000000000000000000000020202222222334455655555444434444545555556667778888888;
		rom_data[190] <= 3840'h7777777777777777777777777777777777777777777777777777777776767776666666666666666666557EEEEEEEC9CEEEEECCCCBAAAABBCBBABAA989A9ABA8778AAA89BCBAAABCCCCCCBCCCCC9999ABAAAAAAAABAAA9ACCCA999AA97898768888CB98ABACABBBCCCBABA999987788BCCA8775578A868AB99989976688767778A97788867765667755AC98AAC9BAABBAA88999A98A889988888758A778656AB988ACECC989A9BAAAA89AAABCCBCCEA8BEEEACCA767777777777777877777776555433332202000000000000000000000000002000022022222333455556555444444444455555555667777888888777777777777777777777777777777777777777777777777777777777777777776767776666666666666666666557EEEEEEEC9CEEEEECCCCBAAAABBCBBABAA989A9ABA8778AAA89BCBAAABCCCCCCBCCCCC9999ABAAAAAAAABAAA9ACCCA999AA97898768888CB98ABACABBBCCCBABA999987788BCCA8775578A868AB99989976688767778A97788867765667755AC98AAC9BAABBAA88999A98A889988888758A778656AB988ACECC989A9BAAAA89AAABCCBCCEA8BEEEACCA767777777777777877777776555433332202000000000000000000000000002000022022222333455556555444444444455555555667777888888;
		rom_data[191] <= 3840'h777777777777777777777777777777777777777777777777777777777767666766666666656665665557CEEEEEEA87BEECECCCBAABBAABCCCA9AA999BA9A98889BB988ACCCBABBCBBCECBBBBCA98899A99ABA998BBAAABECCAA999988ACB999979BB9889BB9AA98ACCCC899888788779BA9A8667888688899778975788778878BA9887778778889976CE879ABABCBBB8CA879BA88A88A9778A9657987889ABA767989BEBAA999ABBA999A9ABBCBCCBABEEEEBECB8767777777777777777766555433322222000000000000000000000000000002020222022233344555555544443444455555555666777787888877777777777777777777777777777777777777777777777777777777777777777767666766666666656665665557CEEEEEEA87BEECECCCBAABBAABCCCA9AA999BA9A98889BB988ACCCBABBCBBCECBBBBCA98899A99ABA998BBAAABECCAA999988ACB999979BB9889BB9AA98ACCCC899888788779BA9A8667888688899778975788778878BA9887778778889976CE879ABABCBBB8CA879BA88A88A9778A9657987889ABA767989BEBAA999ABBA999A9ABBCBCCBABEEEEBECB87677777777777777777665554333222220000000000000000000000000000020202220222333445555555444434444555555556667777878888;
		rom_data[192] <= 3840'h77777777777777777777777777777777777777777777777777777777777676766676666666656665568EEEEEEE975AEECCECBAAAACAABCECB99A9A9AAAAA9989AAA88ABCCCCCCCCCCCCCBABBA9988899999A9988AAAACEEECBA988889CCBA98988A98888A99AA9889BBA88876779A888889B9778888788988787775678889989ABA9877788ACBACCA8AC8579BCBCCBA8BA879AA98977777788866678888BCA886675578ABBBA99BAAA99A99AABBBABCCEEEEEEEEA76777777777777776665555443332220020000000000000000000000000000202020222222234445555555444344445555555566677778888887777777777777777777777777777777777777777777777777777777777777777777676766676666666656665568EEEEEEE975AEECCECBAAAACAABCECB99A9A9AAAAA9989AAA88ABCCCCCCCCCCCCCBABBA9988899999A9988AAAACEEECBA988889CCBA98988A98888A99AA9889BBA88876779A888889B9778888788988787775678889989ABA9877788ACBACCA8AC8579BCBCCBA8BA879AA98977777788866678888BCA886675578ABBBA99BAAA99A99AABBBABCCEEEEEEEEA7677777777777777666555544333222002000000000000000000000000000020202022222223444555555544434444555555556667777888888;
		rom_data[193] <= 3840'h777777777777777777777777777777777777777777777777777777777776777676666666666665557AEEEEEEEA778CECCCCBBBA9BBABCECB99BAAAAA99AAA99AA89ABBBBCCECEEECAABBAAAA999899999A9988888AABCEEEBBA888889AAA8889A888888999BBAA99A9888766789CCCB9877887788888899767996765778ABA889A9888889ABCA89BCB9A9567ABBCCB98A878989C9A877777754788778778A977875677778ABCB999999BA99999BC99ACCEEEECEEC976676777777766555555444333222202000000000000000000000000000000202022022233333455555554444445555555555666777888888877777777777777777777777777777777777777777777777777777777777777777776777676666666666665557AEEEEEEEA778CECCCCBBBA9BBABCECB99BAAAAA99AAA99AA89ABBBBCCECEEECAABBAAAA999899999A9988888AABCEEEBBA888889AAA8889A888888999BBAA99A9888766789CCCB9877887788888899767996765778ABA889A9888889ABCA89BCB9A9567ABBCCB98A878989C9A877777754788778778A977875677778ABCB999999BA99999BC99ACCEEEECEEC9766767777777665555554443332222020000000000000000000000000000002020220222333334555555544444455555555556667778888888;
		rom_data[194] <= 3840'h77777777777777777777777777777777777777777777777777777777777767776777666666665557CEEEEEEEA888EECCCCBABBAAABBCECCBAAABA9AA9888989A99BCCBBCEEEEEECB99ABAB9999899B999BA989988999BEEBA898998777898889C9888999AAABBA89987777778ABCCCCCA876578887778885567755457889999789877778BA898888ABABA66588ACC9988557878BA9999778555799BA976787888989BCB7688AEB8999AAA9999ABECAAAABCECACEEC8666777777775555555444333222220000000000000000000000002022020200220222222233334455555544545555555555566777788888887777777777777777777777777777777777777777777777777777777777777777777767776777666666665557CEEEEEEEA888EECCCCBABBAAABBCECCBAAABA9AA9888989A99BCCBBCEEEEEECB99ABAB9999899B999BA989988999BEEBA898998777898889C9888999AAABBA89987777778ABCCCCCA876578887778885567755457889999789877778BA898888ABABA66588ACC9988557878BA9999778555799BA976787888989BCB7688AEB8999AAA9999ABECAAAABCECACEEC866677777777555555544433322222000000000000000000000000202202020022022222223333445555554454555555555556677778888888;
		rom_data[195] <= 3840'h7777777777777777777777777777777777777777777777777777777777777676766666666655568BEEEEEEEC999CECCCECBABBAAAACCBAAAAAAA99AB988999999ACEBBCEECEEEECB99ABBBAA9888AA99ABA9AA999898BCCA889888877788888ABA88889AA99BA976777788788899A98BCC765799877898877765444789888999766786589889AB9988888575557AB9976457779B98888777777778ACE978978AAC878CEE9977ACB889ABA99AAAABBCEB88C9777ACEB86777676665555544443333222200200000000000000000000022222020200202222222233333444455544454555555555556677778888888777777777777777777777777777777777777777777777777777777777777777777777676766666666655568BEEEEEEEC999CECCCECBABBAAAACCBAAAAAAA99AB988999999ACEBBCEECEEEECB99ABBBAA9888AA99ABA9AA999898BCCA889888877788888ABA88889AA99BA976777788788899A98BCC765799877898877765444789888999766786589889AB9988888575557AB9976457779B98888777777778ACE978978AAC878CEE9977ACB889ABA99AAAABBCEB88C9777ACEB86777676665555544443333222200200000000000000000000022222020200202222222233333444455544454555555555556677778888888;
		rom_data[196] <= 3840'h78777777777777777777777777777777777777777777777777777777777777777776666656557CEEEEEEECC98CBEEECEECBBBAAAABCAA9A99AAA99ABA89AA999AABABCECECCECBAAAABBC99A98889989999BCA998899BCB989878899CCA8789CC8789988888875566789888899AAA889A9667789889CCCCB87566689877ACAA9755887578AAAAABC98875587533688865457778CCB8887778857AC87CE989769CE9348EEE9878CC9899AAAA9AA986BEEB8A745689ACB76676665555554433333232222200000000000000000000022222222220202002020222223333344555554555555555555666777788888887777777778777777777777777777777777777777777777777777777777777777777777777776666656557CEEEEEEECC98CBEEECEECBBBAAAABCAA9A99AAA99ABA89AA999AABABCECECCECBAAAABBC99A98889989999BCA998899BCB989878899CCA8789CC8789988888875566789888899AAA889A9667789889CCCCB87566689877ACAA9755887578AAAAABC98875587533688865457778CCB8887778857AC87CE989769CE9348EEE9878CC9899AAAA9AA986BEEB8A745689ACB7667666555555443333323222220000000000000000000002222222222020200202022222333334455555455555555555566677778888888;
		rom_data[197] <= 3840'h777777777777777777777777777777777777777777777777777777777777777676766665568CEEEEEEEEBB758ABEEEEEECBBAABABBBBBBAA99AA9ABB989AAA9AA99BCECEECBCCA9CBBBA9898988899A989AB988889A9AAAA9988889CB9A888888889A98767875456778999899A9888779A756799ABB988799756768877BB889855788757ABBCB9AAB98547778544554446777779EEB8788788888888BCC898788AC6359EEC866AB988899AA999AA9A9CECA6445998AC966665555554443333322222202000000000000000000002222232222220200202022022233344445555555555555555566677778888888977777777777777777777777777777777777777777777777777777777777777777777777676766665568CEEEEEEEEBB758ABEEEEEECBBAABABBBBBBAA99AA9ABB989AAA9AA99BCECEECBCCA9CBBBA9898988899A989AB988889A9AAAA9988889CB9A888888889A98767875456778999899A9888779A756799ABB988799756768877BB889855788757ABBCB9AAB98547778544554446777779EEB8788788888888BCC898788AC6359EEC866AB988899AA999AA9A9CECA6445998AC9666655555544433333222222020000000000000000000022222322222202002020220222333444455555555555555555666777788888889;
		rom_data[198] <= 3840'h7777777787877777777777777778777777777777777777777777777777777777777666558EEEEA9CEEEEB8559ABEEEEECBBAAAABABBABBAAABBABCCCAAAAABA9AAABCCECECABBAAAAAAA88899899899999888888ABB9ACCBA998889BC9AAA8888999898878866788899AAA88888898A98998778AA9998978997576777BEC788756788889AAAAB899996457778755554577777779CEE9787757899878A99788788BA6348BEE95477898988989AAA99877BEA77748BAABA765555554444333332322202200000000000000000002223333333332222202020202222233344455555555555555666667777788888898777777777777777787877777777777777778777777777777777777777777777777777777777666558EEEEA9CEEEEB8559ABEEEEECBBAAAABABBABBAAABBABCCCAAAAABA9AAABCCECECABBAAAAAAA88899899899999888888ABB9ACCBA998889BC9AAA8888999898878866788899AAA88888898A98998778AA9998978997576777BEC788756788889AAAAB899996457778755554577777779CEE9787757899878A99788788BA6348BEE95477898988989AAA99877BEA77748BAABA765555554444333332322202200000000000000000002223333333332222202020202222233344455555555555555666667777788888898;
		rom_data[199] <= 3840'h77777777778887778777777777787777777777777777777777777777777777777776656AEEEB978EEEEC8755ACEEEEECABBAAAA9AA99BBBBA9ABCCCBBCBBBBBBBBBBCEECCA9BA99999AA988A9899998898898889999AABA99A99999AAA889999BBBBA88AA88678987899AA9788A89AA99BB97789999AAA88877757678ACC777777888899987898878755777787677676778998789CE97788678987667656886767675469BCC77657A9AC9888999999889889CC8ABBCCBA755554444333332322222200020000000000000000022333343433332222202002020222334445555555555555566677777778888899897777777777777777778887778777777777787777777777777777777777777777777777777776656AEEEB978EEEEC8755ACEEEEECABBAAAA9AA99BBBBA9ABCCCBBCBBBBBBBBBBCEECCA9BA99999AA988A9899998898898889999AABA99A99999AAA889999BBBBA88AA88678987899AA9788A89AA99BB97789999AAA88877757678ACC777777888899987898878755777787677676778998789CE97788678987667656886767675469BCC77657A9AC9888999999889889CC8ABBCCBA75555444433333232222220002000000000000000002233334343333222220200202022233444555555555555556667777777888889989;
		rom_data[200] <= 3840'h7777777877877778787777877777877777777777777777777777777777777777776656BEEE9989CEECA988778CEACEECABCAAA999999AA9BBAABCCCBBCBCCECCCCCCCCCBAAABBAB999AAA9999999998888AA778899A988889A9AAAAABBA999889AAA9988987899987886777789BAAA88ABA87787578999777655677778AA87777778765555555555633787777888877767778978AEC97777877755444345787778598657CCC97779B86ACB88999A99BA7558ABACCCCCAB96454433333323223222202200000000000000000222334444545433332222020002022223345555555555565666777777888888899999777777777777777877877778787777877777877777777777777777777777777777777777776656BEEE9989CEECA988778CEACEECABCAAA999999AA9BBAABCCCBBCBCCECCCCCCCCCBAAABBAB999AAA9999999998888AA778899A988889A9AAAAABBA999889AAA9988987899987886777789BAAA88ABA87787578999777655677778AA87777778765555555555633787777888877767778978AEC97777877755444345787778598657CCC97779B86ACB88999A99BA7558ABACCCCCAB96454433333323223222202200000000000000000222334444545433332222020002022223345555555555565666777777888888899999;
		rom_data[201] <= 3840'h7777777777777877777887878778777788888878777777777777777777777777776659EEEB9AAEEEE87788A87AB9EEECCCABAA999989998BECBBBBCCBAABCCCCCEEECEBA99AA9ABA9A999999999A998889B97789AB87777899AAAAAABAAB98777889888888899A9888856777789AA9778976777544675655555576788889A9887788765555444344545777877799977778767757BCC977767575345444568769CA98A9559CCB89AABA559EC9899A89AA987889ABEB9989A7543433222222222222220000000000000000000223344555555444333222220202022233345555556566666667777777888889899999777777777777777777777877777887878778777788888878777777777777777777777777776659EEEB9AAEEEE87788A87AB9EEECCCABAA999989998BECBBBBCCBAABCCCCCEEECEBA99AA9ABA9A999999999A998889B97789AB87777899AAAAAABAAB98777889888888899A9888856777789AA9778976777544675655555576788889A9887788765555444344545777877799977778767757BCC977767575345444568769CA98A9559CCB89AABA559EC9899A89AA987889ABEB9989A7543433222222222222220000000000000000000223344555555444333222220202022233345555556566666667777777888889899999;
		rom_data[202] <= 3840'h777777777877878787877877778787877777788777777777777777777777777776758EEEA89AEEEE988899989BBCEECCCBAA99999988999CCCBCCBBBA9ABBBBBCCCECCB9AA999ABBAA9899A99999999999988887786688889998889997788877888A99999889998898877887788888655556667754554333345675679988AA988788777777656555677658B9779B8777778877667EC978866675467765778669C9C878746CCA8AA99B8448EE98998889CEBA9A9BCC8678A9533333222222222222202200000000000000002233445556555544433322220200022223345555566666666777777777888889999AAA77777777777777777877878787877877778787877777788777777777777777777777777776758EEEA89AEEEE988899989BBCEECCCBAA99999988999CCCBCCBBBA9ABBBBBCCCECCB9AA999ABBAA9899A99999999999988887786688889998889997788877888A99999889998898877887788888655556667754554333345675679988AA988788777777656555677658B9779B8777778877667EC978866675467765778669C9C878746CCA8AA99B8448EE98998889CEBA9A9BCC8678A9533333222222222222202200000000000000002233445556555544433322220200022223345555566666666777777777888889999AAA;
		rom_data[203] <= 3840'h77777878777877787777878878778787878787777777777777777777777777777765BEEC888BEEECA99BCA88BEBBECCEBAAA9999AA989ABBBABCCCCC99ABBBAABCECCBABCB9999AAAA999AB99999999AA98887655668888889876557866689888999AABAA98888788888888888877644455666788755543444576667788899998777667888777878887778BC868A7567768888865BC988867775788876867876888768855CB888888AA5459B98898889ABC9B989CE9688CB7533222222222222202020000000000000000223334556665555554433322202022222333455556666667667777777777888899AAAAA7777777777777878777877787777878878778787878787777777777777777777777777777765BEEC888BEEECA99BCA88BEBBECCEBAAA9999AA989ABBBABCCCCC99ABBBAABCECCBABCB9999AAAA999AB99999999AA98887655668888889876557866689888999AABAA98888788888888888877644455666788755543444576667788899998777667888777878887778BC868A7567768888865BC988867775788876867876888768855CB888888AA5459B98898889ABC9B989CE9688CB7533222222222222202020000000000000000223334556665555554433322202022222333455556666667667777777777888899AAAAA;
		rom_data[204] <= 3840'h77777878888878788878787878787877877788787877777777777777777777777667EEEB988EEECCA99AA87ACBACC9ACCAAAA9A9AA9999ABABCCCABCA9ACAA99BCCAA99CEB9889AA9AA9ACB9AA99999AA998876578898888888765578788998887678778A8887788989888888775555456787757877786677678777657887798755777789A8887777877778B867855777578757648CA88657776776668876776566578868C9789977AB85567569AA98999CC8668AB98CABCA852222222222222202000000000000000002233345556666665554444332222000022334455556666677777777777777788999AAAAA7777777777777878888878788878787878787877877788787877777777777777777777777667EEEB988EEECCA99AA87ACBACC9ACCAAAA9A9AA9999ABABCCCABCA9ACAA99BCCAA99CEB9889AA9AA9ACB9AA99999AA998876578898888888765578788998887678778A8887788989888888775555456787757877786677678777657887798755777789A8887777877778B867855777578757648CA88657776776668876776566578868C9789977AB85567569AA98999CC8668AB98CABCA852222222222222202000000000000000002233345556666665554444332222000022334455556666677777777777777788999AAAAA;
		rom_data[205] <= 3840'h77777777887787878888787877777888778787878777878777777777777777777759EECCB9CEECCCB99A99ACCBCCC79BB999999AAA888999BCBCBBBB9ABA99A9BCB989AEEB888ABA9AAABCB999999ABA8888889A9A98888788778889899988887556655788998878989899888777788888888657668877777778788888888786557998778987777899886556556657776677556667CC8767887665569EEC867877547ACEEEA8998758CB986546878CA999ACB778A88AECBACC7322222222222202002000000000000000223345556667676665554443322020222233345555666777777777766666778889AAAABB7777777777777777887787878888787877777888778787878777878777777777777777777759EECCB9CEECCCB99A99ACCBCCC79BB999999AAA888999BCBCBBBB9ABA99A9BCB989AEEB888ABA9AAABCB999999ABA8888889A9A98888788778889899988887556655788998878989899888777788888888657668877777778788888888786557998778987777899886556556657776677556667CC8767887665569EEC867877547ACEEEA8998758CB986546878CA999ACB778A88AECBACC7322222222222202002000000000000000223345556667676665554443322020222233345555666777777777766666778889AAAABB;
		rom_data[206] <= 3840'h77777787778787878888887778787778787877778787777787777777777777777759ECCB99EECBCB87788BCBBCEE8BCBB99999ACB999A899BCBCBABBBB9989989A9889BCB988AA9AA98899A989ABBBAA99988899A98788878887788899A98888888888888B988877879A988888888988998888789A98987787775798986786667767878755456888ABA87665589875675666677777BB77877757AB97558EE8556AB95569EEC9A99877B899867864589A988AA9999888CBABBCB7322222232222222000000000000000223334455667676776666555433322220222334455556667777777776555566778899AABAB7777777777777787778787878888887778787778787877778787777787777777777777777759ECCB99EECBCB87788BCBBCEE8BCBB99999ACB999A899BCBCBABBBB9989989A9889BCB988AA9AA98899A989ABBBAA99988899A98788878887788899A98888888888888B988877879A988888888988998888789A98987787775798986786667767878755456888ABA87665589875675666677777BB77877757AB97558EE8556AB95569EEC9A99877B899867864589A988AA9999888CBABBCB7322222232222222000000000000000223334455667676776666555433322220222334455556667777777776555566778899AABAB;
		rom_data[207] <= 3840'h7777777778787878888787888787787787878887877787877777777777777777776ACBB989ECCCBA7658ACCBBEEBA899A99999BBA989A999ABBBBAABBCA9AB89999989A999989999A999989ABBCCBABA8A97789A976778777898877789BB7898989B8999CC999898778998788888898899768889AAA8887888855557755667788755668766567877787777788987555855577676698678767767A9878988CE84566855547CECA998855679A88CB9556ABBBA99987888978ACCCB942223232322202000000000000000223345555677777766766655543322202222333455556677777776655555555677899AAABB777777777777777778787878888787888787787787878887877787877777777777777777776ACBB989ECCCBA7658ACCBBEEBA899A99999BBA989A999ABBBBAABBCA9AB89999989A999989999A999989ABBCCBABA8A97789A976778777898877789BB7898989B8999CC999898778998788888898899768889AAA8887888855557755667788755668766567877787777788987555855577676698678767767A9878988CE84566855547CECA998855679A88CB9556ABBBA99987888978ACCCB942223232322202000000000000000223345555677777766766655543322202222333455556677777776655555555677899AAABB;
		rom_data[208] <= 3840'h7777777787877787878788877878777788777787878787777777777777777777776ABBA77CCCBCB7557AAECCCEB9A989AA9899AA9998999999AABACCCCCAAA99889A988998988999A99AA99ABBCBBBA99A888999877788878ABBA987678877888789889AEE999888887897778887888876678889ABB9875567766555456778888777777887888877766677788777555755678875585359856778887679979EE85667655777CEC8789867678888BEB9878ACA989888779888ABABCA4222323222220200000000000002233445556677777777776665544332222222334455556777777665555444445557788AAAAB777777777777777787877787878788877878777788777787878787777777777777777777776ABBA77CCCBCB7557AAECCCEB9A989AA9899AA9998999999AABACCCCCAAA99889A988998988999A99AA99ABBCBBBA99A888999877788878ABBA987678877888789889AEE999888887897778887888876678889ABB9875567766555456778888777777887888877766677788777555755678875585359856778887679979EE85667655777CEC8789867678888BEB9878ACA989888779888ABABCA4222323222220200000000000002233445556677777777776665544332222222334455556777777665555444445557788AAAAB;
		rom_data[209] <= 3840'h77777788787778787888878888778887878778787787778777777777777777777779BB857CCBCB8557BCCCECEEA9AA99A99999A9888889999999ACCCCCB99BAA89AA8889988889899888AABBBBCBCB889988898987788888A9BA9BB9567887787778789CEE99A97788878767887777765689888778A864456766886656677888889BA88987777767777777686567765656888875454337976677888778889CEB77776568987CEA767AB986578669CECA889A99999888ECBA8899CC73232332222020000000000000223344555677777776766776655544332222223344555566766655555433333334557889AABA7777777777777788787778787888878888778887878778787787778777777777777777777779BB857CCBCB8557BCCCECEEA9AA99A99999A9888889999999ACCCCCB99BAA89AA8889988889899888AABBBBCBCB889988898987788888A9BA9BB9567887787778789CEE99A97788878767887777765689888778A864456766886656677888889BA88987777767777777686567765656888875454337976677888778889CEB77776568987CEA767AB986578669CECA889A99999888ECBA8899CC73232332222020000000000000223344555677777776766776655544332222223344555566766655555433333334557889AABA;
		rom_data[210] <= 3840'h7777877777778788887878787878778787787777877887777777777777777777777887557B9AB8558AECCCCBCCB99889A99A9999889998998999ACCCCBA89A9899AA88899887899998889ABBCCBBB8589899878887787789979989B9778987777888889CECABBA77888666789768998778989886555544567777875887777776689CCAA977775677887876775567787777788877677635BC8656789898779BA8775787789A78CE9779CCB85797359BEEEA7789AAA999CAA9888AA9853232322220200000000000222334455567777777776776676655544333322233345555666655554433333222334567899AAA777777777777877777778788887878787878778787787777877887777777777777777777777887557B9AB8558AECCCCBCCB99889A99A9999889998998999ACCCCBA89A9899AA88899887899998889ABBCCBBB8589899878887787789979989B9778987777888889CECABBA77888666789768998778989886555544567777875887777776689CCAA977775677887876775567787777788877677635BC8656789898779BA8775787789A78CE9779CCB85797359BEEEA7789AAA999CAA9888AA9853232322220200000000000222334455567777777776776676655544333322233345555666655554433333222334567899AAA;
		rom_data[211] <= 3840'h77777878787878888888788887877878787878877787787877777777777777777768756897887558BCCCCCCB9AA9778999AA9999988999999988BCBBCCA999889AB9888898788999988899AAA8888768A89A875788777799889A9988778887778A989988AA99B9778887678987799AA9AA978887554446676677555997787776558CB898788778889878877557887777665787789AC944ACA6456889987778656556998889878EC8878CEB88A843589CEE968ABAAA99878789BCC88732232222020000000000022233445556677777777777777766655543332232334445555555554433322222222334577899AA7777777777777878787878888888788887877878787878877787787877777777777777777768756897887558BCCCCCCB9AA9778999AA9999988999999988BCBBCCA999889AB9888898788999988899AAA8888768A89A875788777799889A9988778887778A989988AA99B9778887678987799AA9AA978887554446676677555997787776558CB898788778889878877557887777665787789AC944ACA6456889987778656556998889878EC8878CEB88A843589CEE968ABAAA99878789BCC88732232222020000000000022233445556677777777777777766655543332232334445555555554433322222222334577899AA;
		rom_data[212] <= 3840'h7778777787777887887887888887877778878778787877777777777777777777778A78CE9765459AACBECBCB878778999A999999888889A9AA88BCCCCCAAAAA99A98888888888898888888875445688888998657886899BAABCBB9876788887799999A988876775688887998888987789BB85677778767766675557877787798747CC877788899789888887667CB6577556888778AA8548C955556876787655455658879B9878BC97657B989A7434668CEECCBCA9A9867A9ACCECBA84223222202000000000222233445556667777777777777767766555443332323344555555444333222202000223446778899777777777778777787777887887887888887877778878778787877777777777777777777778A78CE9765459AACBECBCB878778999A999999888889A9AA88BCCCCCAAAAA99A98888888888898888888875445688888998657886899BAABCBB9876788887799999A988876775688887998888987789BB85677778767766675557877787798747CC877788899789888887667CB6577556888778AA8548C955556876787655455658879B9878BC97657B989A7434668CEECCBCA9A9867A9ACCECBA84223222202000000000222233445556667777777777777767766555443332323344555555444333222202000223446778899;
		rom_data[213] <= 3840'h7777787877878788888888878878888887787877777777777777777777777777779CCCEE76556899AAECCB9A97777AA9A988999989888998999ABCCCCBBCABA99988788888888888887888654444688779BA878A88579AAA9ACCA98757887777899AA98998755557889888888888867878A86666789778756655668766788888767AB8877779A8776899765545A96775556887748A99658CA5654455555665544675775799777AB98854788987533468ACCCB99A99A998BCCAAABBB95232222220000000002223333445566777777777767777677766555543332333343445444433322202000002223345577888767777777777787877878788888888878878888887787877777777777777777777777777779CCCEE76556899AAECCB9A97777AA9A988999989888998999ABCCCCBBCABA99988788888888888887888654444688779BA878A88579AAA9ACCA98757887777899AA98998755557889888888888867878A86666789778756655668766788888767AB8877779A8776899765545A96775556887748A99658CA5654455555665544675775799777AB98854788987533468ACCCB99A99A998BCCAAABBB95232222220000000002223333445566777777777767777677766555543332333343445444433322202000002223345577888;
		rom_data[214] <= 3840'h777777787787778888787887888878888878777887777877777777777777777777BCCEEC555789BBBEEEA89BB877ABAAA988898888888999989ACCCCBABCCBBB999878888888889887887655555788889AAA877877668A9989BB987547887787888888887887778877888898888777888789767889877767676577655657998678ACB89877788567678854555555567654678865598877ABA55543334445554457876555788879B988855689776533578AB9A8789A9998ACCCA88ACC842222202020000002223334455566777777777777777777777665554433323333444444333222200000000002233555677877777777777777787787778888787887888878888878777887777877777777777777777777BCCEEC555789BBBEEEA89BB877ABAAA988898888888999989ACCCCBABCCBBB999878888888889887887655555788889AAA877877668A9989BB987547887787888888887887778877888898888777888789767889877767676577655657998678ACB89877788567678854555555567654678865598877ABA55543334445554457876555788879B988855689776533578AB9A8789A9998ACCCA88ACC8422222020200000022233344555667777777777777777777776655544333233334444443332222000000000022335556778;
		rom_data[215] <= 3840'h777777787878787888888887888888787887888877878777777777777777777778EEEEEB78ACABCBCEEC989ABB98BCA888988999988CCB98988ABABCCBBCBBBA999888789988889777877777888998899A9986788777789877998753588778888888998889888788789A9998767788A988778778888877877556888667668986757AA88767555678767545777755675433578855557878A67577433222334345777885345788789977975668CB7333357787677678AA988BBBB88ACEEA4222020200000022233344555667677777777777777777777766555443333333334333323220000000000222223455556767777777777777787878787888888887888888787887888877878777777777777777777778EEEEEB78ACABCBCEEC989ABB98BCA888988999988CCB98988ABABCCBBCBBBA999888789988889777877777888998899A9986788777789877998753588778888888998889888788789A9998767788A988778778888877877556888667668986757AA88767555678767545777755675433578855557878A67577433222334345777885345788789977975668CB7333357787677678AA988BBBB88ACEEA42220202000000222333445556676777777777777777777777665554433333333343333232200000000002222234555567;
		rom_data[216] <= 3840'h77777778787878888788888887878787887878787878777777777777777777778EEEECACCCEC89ABEEE8899ABAA9CB988888999889ACA88A989AAABCCCBBBBCBA98888888A988888887788887799878877677579887678877689853478778AAA8678AA88AA98888767ACCA97555789A98898887777877687665578755755567557778788777679887555578787777655547756765357786345865545332233687535875345788987778657768AE95323555555779ABA99999ABAABABEE730220000000022233444555567777777777777777777777776655544433333333333322222000000000000022234455557777777777777778787878888788888887878787887878787878777777777777777777778EEEECACCCEC89ABEEE8899ABAA9CB988888999889ACA88A989AAABCCCBBBBCBA98888888A988888887788887799878877677579887678877689853478778AAA8678AA88AA98888767ACCA97555789A98898887777877687665578755755567557778788777679887555578787777655547756765357786345865545332233687535875345788987778657768AE95323555555779ABA99999ABAABABEE73022000000002223344455556777777777777777777777777665554443333333333332222200000000000002223445555;
		rom_data[217] <= 3840'h7777777878887878888888888888888887787877778777777777777777777777AEEEEACEEBCB89ACEE878989BAAACA888888998889AA879BA89A99BCCCBAAAABA88889889998887788778887666777885565558998755777777753357878ABA8758AB889AA77888875789BB7554688988AA887777776788756654454576755545887778878778A9776555788988865565665588785456642456556567554467775345655345799775556577657BEB633343444589CCC99999A9AA8778A94020020000222333444555666777777777777777777777777776555444333333333222200000000000020222223334445777777777777777878887878888888888888888887787877778777777777777777777777AEEEEACEEBCB89ACEE878989BAAACA888888998889AA879BA89A99BCCCBAAAABA88889889998887788778887666777885565558998755777777753357878ABA8758AB889AA77888875789BB7554688988AA887777776788756654454576755545887778878778A9776555788988865565665588785456642456556567554467775345655345799775556577657BEB633343444589CCC99999A9AA8778A94020020000222333444555666777777777777777777777777776555444333333333222200000000000020222223334445;
		rom_data[218] <= 3840'h7777777877788888788888888787888878787878887877777777777777777778EEEEBACEC9BB8ACEE9889979B9AAA988998888888AA688AA989988ABBBAAAA999889999999888888887788777765779A55555789A875455555544458888899875589A8778757AA8886556997674567778A9996557876567555764455677877567888788888878988776657777865557777557987864455336565566775656887986555565345688655565575557AEB733333457878BCAB99998887788995202000000222333455556677777777777777777777777777776655544433333232222000000000000000002222233344677777777777777877788888788888888787888878787878887877777777777777777778EEEEBACEC9BB8ACEE9889979B9AAA988998888888AA688AA989988ABBBAAAA999889999999888888887788777765779A55555789A875455555544458888899875589A8778757AA8886556997674567778A9996557876567555764455677877567888788888878988776657777865557777557987864455336565566775656887986555565345688655565575557AEB733333457878BCAB99998887788995202000000222333455556677777777777777777777777777776655544433333232222000000000000000002222233344;
		rom_data[219] <= 3840'h777777777787888888788888888887878888878777777777777777777777767BEEEB98BC8ACA9AEE98A99878B8989889888888889B959A88888888BBBAAABA9899899998988889A988788877777678A97557788998764444434556999A887776568898655558988898556765896445568988964588754433467755687777788888888988998778987787577555555687877899887743543487785555455567768876756765444555555655665558BEB5322348BA77ABAAA89887679CAAA722000000222333455556777777777777777777777777777777766555443333222220000000000000000202202222333377777777777777777787888888788888888887878888878777777777777777777777767BEEEB98BC8ACA9AEE98A99878B8989889888888889B959A88888888BBBAAABA9899899998988889A988788877777678A97557788998764444434556999A887776568898655558988898556765896445568988964588754433467755687777788888888988998778987787577555555687877899887743543487785555455567768876756765444555555655665558BEB5322348BA77ABAAA89887679CAAA7220000002223334555567777777777777777777777777777777665554433332222200000000000000002022022223333;
		rom_data[220] <= 3840'h777777778788787888878888878887878787888887878777777777777777758EEEC878AB9CC99EEC89B98888A999998888888888BC77997888888ABAAAAAAA988999A88888999AA88888987887779A9875677778778864444577777789777775688899755778777898878755888533567787854588765444577556677888778988768878875557886776677655666776788AA8787643323577775444475576555676557757544334434665678558ACA7422258ABCA9A99A989876ACCCBA720200002022344555667777777777777777777777777777777776555444333322020000000000000000000022222222377677777777777778788787888878888878887878787888887878777777777777777758EEEC878AB9CC99EEC89B98888A999998888888888BC77997888888ABAAAAAAA988999A88888999AA88888987887779A9875677778778864444577777789777775688899755778777898878755888533567787854588765444577556677888778988768878875557886776677655666776788AA8787643323577775444475576555676557757544334434665678558ACA7422258ABCA9A99A989876ACCCBA7202000020223445556677777777777777777777777777777777765554443333220200000000000000000000222222223;
		rom_data[221] <= 3840'h777777787878888878888888888887878887878878787777777777777777769CEEB989BCECA8AEECBBB987899999B98888888988CA6A87788899ABAA99A999989A89A9998899988889A876899889AA8777667765788888777988754357799977897899778987888889A98777658753455555655587777666777777556888768A97567767543567777566765777777778889A964655433236575443435A6565455678547756545543223775588658898565335747988CA99999987BECCB9632000020223345556777777777777777777777777777777777777655544333222200000000000000000002222222223376777777777777787878888878888888888887878887878878787777777777777777769CEEB989BCECA8AEECBBB987899999B98888888988CA6A87788899ABAA99A999989A89A9998899988889A876899889AA8777667765788888777988754357799977897899778987888889A98777658753455555655587777666777777556888768A97567767543567777566765777777778889A964655433236575443435A6565455678547756545543223775588658898565335747988CA99999987BECCB96320000202233455567777777777777777777777777777777777776555443332222000000000000000000022222222233;
		rom_data[222] <= 3840'h777777777778787888788888788788878788887878787877777777777777777BCCA978CCCA789CECCBA987799889988888888A8BB77A88987899998999999899A99889B989AA8889998657876888876566677755778889877778755557799777767999987788A97667877787667774334543335677665567777566778888754687678768667776689899867875777899888854576433333555567655576775457588776565666888655665787658765556577645547CA998999888B9899832202002223445566777777777777777777777777777777777777655544332222000000000000000000000202222232366777777777777777778787888788888788788878788887878787877777777777777777BCCA978CCCA789CECCBA987799889988888888A8BB77A88987899998999999899A99889B989AA8889998657876888876566677755778889877778755557799777767999987788A97667877787667774334543335677665567777566778888754687678768667776689899867875777899888854576433333555567655576775457588776565666888655665787658765556577645547CA998999888B98998322020022234455667777777777777777777777777777777777776555443322220000000000000000000002022222323;
		rom_data[223] <= 3840'h7777777878878888888888788888888888878888878787877777777777778658CCA77A9BE889CECAA9AA8889888998888898987CA57989988998899A889A9889999989BBAAA98888987778899988988888555577788778766778777667788888878AAC9777888988767778987567754333333466666656555654566899888755555785577755787798897457757767886555545654323357655577766456655555766778A756569A755555456768756556787767768C8998888998865589520200202334455677777777777777777777777777777777777776555443332200000000000000000000002222233233677777777777777878878888888888788888888888878888878787877777777777778658CCA77A9BE889CECAA9AA8889888998888898987CA57989988998899A889A9889999989BBAAA98888987778899988988888555577788778766778777667788888878AAC9777888988767778987567754333333466666656555654566899888755555785577755787798897457757767886555545654323357655577766456655555766778A756569A755555456768756556787767768C8998888998865589520200202334455677777777777777777777777777777777777776555443332200000000000000000000002222233233;
		rom_data[224] <= 3840'h7777777777787778888788888888888888888787877778787777777777767779BA859BBC989BECBCA999878988998888889996AC878888779A88A98988999888888899BEBA99888887789A998889A998AA8875788888887775787888778898888799A97677987888876778975566677532223577777656643334777789878877767776776766778787888655546765653334444442245566545455555445565565655559CA57547A9775773235678776567768856876798888889875547B732000222344556777777777777777777777777777777777777777555443322220000000000000000000020222233333666777777777777777787778888788888888888888888787877778787777777777767779BA859BBC989BECBCA999878988998888889996AC878888779A88A98988999888888899BEBA99888887789A998889A998AA8875788888887775787888778898888799A97677987888876778975566677532223577777656643334777789878877767776776766778787888655546765653334444442245566545455555445565565655559CA57547A9775773235678776567768856876798888889875547B732000222344556777777777777777777777777777777777777777555443322220000000000000000000020222233333;
		rom_data[225] <= 3840'h7777777778777888888888888888888888888888878787777777777777669C9888569ABCA78AECBBA975689888988888899A99E858A8888899899888ABB88998889889CECA9888888778888878ABA88788888778888899888677788988988888877675577575689886787755575767A8654577888776776543357765675588777888777677775598A8669B97456776533323323332355578876543455545676785435557BB545668B986765322468986568766867987889A88888888755BB52020223445556777777777777777777777777777777777777777655543322200000000000000000000022223333434667777777777777778777888888888888888888888888888878787777777777777669C9888569ABCA78AECBBA975689888988888899A99E858A8888899899888ABB88998889889CECA9888888778888878ABA88788888778888899888677788988988888877675577575689886787755575767A8654577888776776543357765675588777888777677775598A8669B97456776533323323332355578876543455545676785435557BB545668B986765322468986568766867987889A88888888755BB52020223445556777777777777777777777777777777777777777655543322200000000000000000000022223333434;
		rom_data[226] <= 3840'h77777777777777888888888888888888888878878787878877777777777BCB98656988BCA789CBAA985468888888888889BB8CC878988877888888889A989A98988889BBAA988788887776776898655556788976756678998777765678887888865554588756888877888655775657A98788888877757555555657765556898878A878776576579887558CC9577577657545543332466557878854555554359B85535445885447779A875577422355554586545568B877AA87888999966AB720222334555677777777777777777777777777777777777777766555443322200000000000000000000223333444456667777777777777777777888888888888888888888878878787878877777777777BCB98656988BCA789CBAA985468888888888889BB8CC878988877888888889A989A98988889BBAA988788887776776898655556788976756678998777765678887888865554588756888877888655775657A98788888877757555555657765556898878A878776576579887558CC9577577657545543332466557878854555554359B85535445885447779A875577422355554586545568B877AA87888999966AB72022233455567777777777777777777777777777777777777776655544332220000000000000000000022333344445;
		rom_data[227] <= 3840'h7777777777887878788888888888888888878878877878777777777777BCCCA6559B99BA87BB9AAA95457888888888889ACB9CB9998886578878788788889A9999878998898887778877544455654344545567777776677777765544578777888877678AA858888888977777777557AA8787677778755557765556787567878868B87898667768867775688978646778877775555457765755787555556645AC6575533455465556799674586323343345777635689767B9778888988778974222334555567777777777777777777777777777777777777777665554332202000000000000000000222334444555677777777777777777887878788888888888888888878878877878777777777777BCCCA6559B99BA87BB9AAA95457888888888889ACB9CB9998886578878788788889A9999878998898887778877544455654344545567777776677777765544578777888877678AA858888888977777777557AA8787677778755557765556787567878868B87898667768867775688978646778877775555457765755787555556645AC6575533455465556799674586323343345777635689767B9778888988778974222334555567777777777777777777777777777777777777777665554332202000000000000000000222334444555;
		rom_data[228] <= 3840'h7777777787788887878888888888888888888887878787787777777779CABEB668BACA8779EC88A974478988988888889CC9BBA9999975589877788788889A9AA9889A88898888778887533333344444432334588ACA75545676555567777778898889BCA778888888755776787757AB9765557888755557655557677778757758CA88A878878888988876586A745767757765677677767754457756777887BB5557542333475435578575677644555358878757865577B9888888877888887323345556677777777777777777777777777777777777777777665544322200000000000000000002233344455555666777777777777787788887878888888888888888888887878787787777777779CABEB668BACA8779EC88A974478988988888889CC9BBA9999975589877788788889A9AA9889A88898888778887533333344444432334588ACA75545676555567777778898889BCA778888888755776787757AB9765557888755557655557677778757758CA88A878878888988876586A745767757765677677767754457756777887BB5557542333475435578575677644555358878757865577B9888888877888887323345556677777777777777777777777777777777777777777665544322200000000000000000002233344455555;
		rom_data[229] <= 3840'h777777777787888888888888888878888888878887787777777777779CC9EE989CB9C9558CCB66985468898898888888AEBBBA8899988778988767778888899A98889888898888877778765544333344332333578ACC8544567777787777777898778ABC95888888865565656777779B9876557887545555447877777778968868EEC998777789999A988865687557776667777776555565433487578777889B5555754454686544556565787755557777877678864597AA998888888AA88AB53345555677777777777777777777777777777777777777777777655433222000000000000000002223344455556667777777777777777787888888888888888878888888878887787777777777779CC9EE989CB9C9558CCB66985468898898888888AEBBBA8899988778988767778888899A98889888898888877778765544333344332333578ACC8544567777787777777898778ABC95888888865565656777779B9876557887545555447877777778968868EEC998777789999A988865687557776667777776555565433487578777889B5555754454686544556565787755557777877678864597AA998888888AA88AB533455556777777777777777777777777777777777777777777776554332220000000000000000022233444555566;
		rom_data[230] <= 3840'h7777777777887878878888887888878888888888887887877777778ACC9BCC99CC8AC857CCAC65754798888898988988ABAB998889878878887767887788888988888888898899877777888776322332335566787898765787777568889877788777678865788888877875555557869A9987755565345555556765788678878879EEC88654577888ABA88875554357788867888754335575333576567787779B55555655588866554555755787555578877874666776B788CB878889ABCA8BC843455667777777777777777777777777777777777777777777776555332202000000000000000022234455555666676777777777777777887878878888887888878888888888887887877777778ACC9BCC99CC8AC857CCAC65754798888898988988ABAB998889878878887767887788888988888888898899877777888776322332335566787898765787777568889877788777678865788888877875555557869A9987755565345555556765788678878879EEC88654577888ABA88875554357788867888754335575333576567787779B55555655588866554555755787555578877874666776B788CB878889ABCA8BC843455667777777777777777777777777777777777777777777776555332202000000000000000022234455555666;
		rom_data[231] <= 3840'h7777777877787878888888888788888888888887878877778777779CBA7ACA77A96BCAACEBBC75556997889AA8888888AB888568778777898777787777888888778988877777898778767777776433356765776778876789888777888987677777787555557888878888855576877779A987767676577355555778787777778789ABB875765578889AA887798533565787755555323577556776545678988789566545554697555557655557B956787678555787544477878A88788877BC8AB754556777777777777777777777777777777777777777777777776554433220000000000000002223334555566767666777777777777877787878888888888788888888888887878877778777779CBA7ACA77A96BCAACEBBC75556997889AA8888888AB888568778777898777787777888888778988877777898778767777776433356765776778876789888777888987677777787555557888878888855576877779A987767676577355555778787777778789ABB875765578889AA887798533565787755555323577556776545678988789566545554697555557655557B956787678555787544477878A88788877BC8AB754556777777777777777777777777777777777777777777777776554433220000000000000002223334555566767;
		rom_data[232] <= 3840'h777777777878788778788878788787888888888888888787877778BC77689889978CAAECBBCC64456768988998888878A986545557777897777778777778898888887777788888888887788777765677777555677788889898777787775456788878656778888877889A975688765578998877777755435665688889856886578779CA8776435788889878885434677877766544455665556755544568A98777556555775457757877765766875888646755358A9755555675688988758EA8987555677777777777777777777777777777777777777777777777755443320200000000000000222344455556677766677777777777777878788778788878788787888888888888888787877778BC77689889978CAAECBBCC64456768988998888878A986545557777897777778777778898888887777788888888887788777765677777555677788889898777787775456788878656778888877889A975688765578998877777755435665688889856886578779CA8776435788889878885434677877766544455665556755544568A98777556555775457757877765766875888646755358A9755555675688988758EA89875556777777777777777777777777777777777777777777777777554433202000000000000002223444555566777;
		rom_data[233] <= 3840'h777777778777887788888877888888888888887878787777777779C95698658CA8BB9ACC9CCC534787889899888888899897744457788998787887778778888888877787777888888877887777777777668766777677765556765565554577788776678778778876567A976788577677788877777765457665677877657877777768BB857653467778987886433478755657875555555556985555455687777655755565444575556775555676588754585766799876567777798988857CC8689756777778877777777777777778777777777777877777777777665443222000000000000002223345555667777766677777777777778777887788888877888888888888887878787777777779C95698658CA8BB9ACC9CCC534787889899888888899897744457788998787887778778888888877787777888888877887777777777668766777677765556765565554577788776678778778876567A976788577677788877777765457665677877657877777768BB857653467778987886433478755657875555555556985555455687777655755565444575556775555676588754585766799876567777798988857CC86897567777788777777777777777787777777777778777777777776654432220000000000000022233455556677777;
		rom_data[234] <= 3840'h77777777778778888888888877888888888888878887878787777BC768B977CEEBC88BCA8CCB988899889998888888888AA987555679B9999878877777888888888777877777788877788756777765557887578887655445677655544447887878767887566788877558A757875787777678887777765566543455554478777877668855785435556788776542457874578887655555544798655554246677654555567864557555775455556767975468558878887769BA98788888A87BC858A86777777877778878787777787778777777778777777777777776544332220000000000022223445556666777776666777777777777778778888888888877888888888888878887878787777BC768B977CEEBC88BCA8CCB988899889998888888888AA987555679B9999878877777888888888777877777788877788756777765557887578887655445677655544447887878767887566788877558A757875787777678887777765566543455554478777877668855785435556788776542457874578887655555544798655554246677654555567864557555775455556767975468558878887769BA98788888A87BC858A8677777787777887878777778777877777777877777777777777654433222000000000002222344555666677777;
		rom_data[235] <= 3840'h77777777778787888878878788888878888888888878787877879B879CECACEECACBACA778ACEE98AA8888888888888988888777557CEA99877877777777787888777787777567855578755677766558876556667777555788767754346787778887888776777878875675655577787776578987677555555433334325787776677665566665434455777664335577656787777645776556776545542355555435558779A6675677863355556556556666557776776657CBB9788888BB88AA78A87777888878888777778878887878778788877888887878887776554322000000000000222233455556777777776667777777777777778787888878878788888878888888888878787877879B879CECACEECACBACA778ACEE98AA8888888888888988888777557CEA99877877777777787888777787777567855578755677766558876556667777555788767754346787778887888776777878875675655577787776578987677555555433334325787776677665566665434455777664335577656787777645776556776545542355555435558779A6675677863355556556556666557776776657CBB9788888BB88AA78A8777788887888877777887888787877878887788888787888777655432200000000000022223345555677777777;
		rom_data[236] <= 3840'h77777777777777878788888888787888787887878787777787779A88CEEBCEEB89CCCE8579AEEA57A97888889888788987777788768CCA97678778787778777888777777887556644578655666666778855565545778767887678875578777788887788887676778874546775586656776557995576545545532232246767776577655885567533444577653355655457655567755578777655545543234554344668867B75856887554675676575577558875877776558ABA9877789B877988887888888887888788887787888787787887788777778888787776554322202000000022223333555567677776666666777777777777777777878788888888787888787887878787777787779A88CEEBCEEB89CCCE8579AEEA57A97888889888788987777788768CCA97678778787778777888777777887556644578655666666778855565545778767887678875578777788887788887676778874546775586656776557995576545545532232246767776577655885567533444577653355655457655567755578777655545543234554344668867B75856887554675676575577558875877776558ABA9877789B87798888788888888788878888778788878778788778877777888878777655432220200000002222333355556767777666;
		rom_data[237] <= 3840'h7777777787878877788888787878787887878878887777778777998BEEA8AEC97ACCEC868CCEA55798899889888878889AA7789988ABB9867987778887777787787777888877764456776676666555767656775556777788855778888888777888877789876657777655578998775457776557645777553555533334776577775677678755676443344565332467544577556577654577875455555453224443457757778756677656977757A9887876569A549B87777678888777788998777787788888888888888888887788888887887888888888878788777655433200000202222223333555566777776566666777777777777787878877788888787878787887878878887777778777998BEEA8AEC97ACCEC868CCEA55798899889888878889AA7789988ABB9867987778887777787787777888877764456776676666555767656775556777788855778888888777888877789876657777655578998775457776557645777553555533334776577775677678755676443344565332467544577556577654577875455555453224443457757778756677656977757A9887876569A549B87777678888777788998777787788888888888888888887788888887887888888888878788777655433200000202222223333555566777776566;
		rom_data[238] <= 3840'h7777777778777778878788888787878788888777887877777777889CEC87CC978BBCEB8889EC77899788989888888878EE9567877AA888888887777788877887787777898888754567557777776567788856777788756777745788899887778889877887777568766787877887776577657645446877555655555656876788887776676665557544333443323477776688776577554456555435654553223343458745676454575457775578885558766556548A75765455557777888899887788788888888888888888888888888888888888888888888888887755432220202022222333344555566777665655666677777777777778777778878788888787878788888777887877777777889CEC87CC978BBCEB8889EC77899788989888888878EE9567877AA888888887777788877887787777898888754567557777776567788856777788756777745788899887778889877887777568766787877887776577657645446877555655555656876788887776676665557544333443323477776688776577554456555435654553223343458745676454575457775578885558766556548A75765455557777888899887788788888888888888888888888888888888888888888888888887755432220202022222333344555566777665655;
		rom_data[239] <= 3840'h7777777777777887888877888888887877777887777777777777899AEA88AB867BAEC8888BEA8779A78988887888877AEA6778778888788887777787788878887877778988876557875687778866788887677776777655565367777AB866678999855566677778766888777776675555456755567765555555675556777888998755677886558753323333224555665685565555545554456436654455333334446554555435666567787588655438876433557865665445557788888888888787788888888888888888888888888888888888888888888888887755433200002022223333444555566666655555666777777777777777777887888877888888887877777887777777777777899AEA88AB867BAEC8888BEA8779A78988887888877AEA6778778888788887777787788878887877778988876557875687778866788887677776777655565367777AB866678999855566677778766888777776675555456755567765555555675556777888998755677886558753323333224555665685565555545554456436654455333334446554555435666567787588655438876433557865665445557788888888888787788888888888888888888888888888888888888888888888887755433200002022223333444555566666655555;
		rom_data[240] <= 3840'h77777777777877778888787777887787778777787878777777788A98B87787558ABCA888AEC98677778988887788777BB56987777888567877777788888888787887787877876789888887788657898787665443456765553476558CB8776789998577777788888668877777555444555566777877555777544545576668998885577789A74586544554323355556555455555555555533464455545675654457777555433477677776A65555543466754546558755665434558988888888777767888888888888888888888888888888888888888888888888877654322220202222333444445555556565555556666677777777777777877778888787777887787778777787878777777788A98B87787558ABCA888AEC98677778988887788777BB56987777888567877777788888888787887787877876789888887788657898787665443456765553476558CB8776789998577777788888668877777555444555566777877555777544545576668998885577789A74586544554323355556555455555555555533464455545675654457777555433477677776A6555554346675454655875566543455898888888877776788888888888888888888888888888888888888888888888887765432222020222233344444555555656555555;
		rom_data[241] <= 3840'h7777777777777778878887878877877787777787777777777779AA9885677547AACB9977BE975577788988988887779C95797788888978885677788878788877778877788887789877898776756767778554433455577653467765797576789AB975677777756765687788777645556776578756754455654454455556789B7655677668B8567544775544465656765556777767886543234445544568765345567555543347665577486753345535568876755787458755457898888788886676788888888888888888888888888888888888888888888888887775543220202223333344455555555555555555666767777777777777777778878887878877877787777787777777777779AA9885677547AACB9977BE975577788988988887779C95797788888978885677788878788877778877788887789877898776756767778554433455577653467765797576789AB975677777756765687788777645556776578756754455654454455556789B7655677668B8567544775544465656765556777767886543234445544568765345567555543347665577486753345535568876755787458755457898888788886676788888888888888888888888888888888888888888888888887775543220202223333344455555555555555555;
		rom_data[242] <= 3840'h777777777777787788878878777878787777777777777777778BB887558A745BCACA8768CB86458888988988777777AC87998878888A989777877788888888877778777888789986667887555665445776543457566777766777766755756889A755677775555544677886567757778865777754433543333455665457778975557775557557765577655677565455465776777666555544533455555655544335544555555556655556554456576345775645557974788755699878877898778778888888888888888888888888888888888888888888888888876554322202222333444445445444555544444466676767777777777777787788878878777878787777777777777777778BB887558A745BCACA8768CB86458888988988777777AC87998878888A989777877788888888877778777888789986667887555665445776543457566777766777766755756889A7556777755555446778865677577788657777544335433334556654577789755577755575577655776556775654554657767776665555445334555556555443355445555555566555565544565763457756455579747887556998788778987787788888888888888888888888888888888888888888888888888765543222022223334444454454445555444444;
		rom_data[243] <= 3840'h777777777777777777877877877777777777777787777777778CB88878AA659CB9CA8769E875479988888987777778BB88B98876789988788888777888887887777777778888876667788755676545577543478757777677777777777775578886447766566654567657545565587885556887553346544445655655676556545777755555677757765557885665444677556555555555556545554543344542345545556555555554434567655684557757565569A54789B979BB888878A9777789888888888888888888888888888888888888888888888888877554332202223334445555454444444434343466676777777777777777777777877877877777777777777787777777778CB88878AA659CB9CA8769E875479988888987777778BB88B98876789988788888777888887887777777778888876667788755676545577543478757777677777777777775578886447766566654567657545565587885556887553346544445655655676556545777755555677757765557885665444677556555555555556545554543344542345545556555555554434567655684557757565569A54789B979BB888878A97777898888888888888888888888888888888888888888888888888775543322022233344455554544444444343434;
		rom_data[244] <= 3840'h777777777777777777787777777777777777777777777777779CB88BB88878CCA8998778975459A989888877777879B988A8876678877657888777787788AA88877877777776556888898777888656777544687668997677765678999876567775357875568877787544355544678754455787555457755577655557887544447875556677677667565556776777566787566555556555545556555553344543345555556445554565443775555575557747654457854468ACB9998888879A8757AA888888888888888888888888888888888888888888888888877654432222223334445555443433333333333366666767777777777777777777787777777777777777777777777777779CB88BB88878CCA8998778975459A989888877777879B988A8876678877657888777787788AA88877877777776556888898777888656777544687668997677765678999876567775357875568877787544355544678754455787555457755577655557887544447875556677677667565556776777566787566555556555545556555553344543345555556445554565443775555575557747654457854468ACB9998888879A8757AA8888888888888888888888888888888888888888888888888776544322222233344455554434333333333333;
		rom_data[245] <= 3840'h77777777777777777778777777777777777777777777777778AB999AA7998ABBC8787788665479988988887777887CB8877777778875544567777788788BEB98888887777775556788988787787777777656767787886577656678AA985555566446787667898A9876554675457665556655655565656555566555579986555589756876886787654566654567777877755776556675555445556766544555454335544555455557774557545654345544454553455445557BEA656888878A85579888888888888888888888888888888888888888888888888888765543322223334455555444433333233333336667677777777777777777777778777777777777777777777777777778AB999AA7998ABBC8787788665479988988887777887CB8877777778875544567777788788BEB98888887777775556788988787787777777656767787886577656678AA985555566446787667898A9876554675457665556655655565656555566555579986555589756876886787654566654567777877755776556675555445556766544555454335544555455557774557545654345544454553455445557BEA656888878A8557988888888888888888888888888888888888888888888888888876554332222333445555544443333323333333;
		rom_data[246] <= 3840'h77777777777777777777778778777777777777777777777789A89B988CC99AACB8575776554589889988888787877B98766777788753553567777888888BEB8888888777777776556776766555566577777667756554457756656899864555455356565576788CB8888657656786556887555457755443554354556688887777887688658877775445677545777588544468974557755555455455555557765553235435555555777745555578433564234446643343455679CA545788779995677788898888888888888888888888888888888888888888888888776543332223344455555544433322222223336666766777777777777777777777778778777777777777777777777789A89B988CC99AACB8575776554589889988888787877B98766777788753553567777888888BEB8888888777777776556776766555566577777667756554457756656899864555455356565576788CB8888657656786556887555457755443554354556688887777887688658877775445677545777588544468974557755555455455555557765553235435555555777745555578433564234446643343455679CA54578877999567778889888888888888888888888888888888888888888888888877654333222334445555554443332222222333;
		rom_data[247] <= 3840'h77777777777777777777777777777777777777777777777799789A989B89CECCB95657755558988888888877777787777876677775557745677888888888A878777888777777776555545555445665678767776444445788775458CB755553444366544675567898997554457875676765455588654545554445577777787787665578557657766666554458776677444577655568775555555543455556776554334565555555666654435569657687535355553344356557AA755778778898887678898888989888888888888888888888888888888888888888876554332323344455555544333222222232336666677777777777777777777777777777777777777777777777777799789A989B89CECCB95657755558988888888877777787777876677775557745677888888888A878777888777777776555545555445665678767776444445788775458CB755553444366544675567898997554457875676765455588654545554445577777787787665578557657766666554458776677444577655568775555555543455556776554334565555555666654435569657687535355553344356557AA75577877889888767889888898988888888888888888888888888888888888888887655433232334445555554433322222223233;
		rom_data[248] <= 3840'h777777777777777777777777777777777777777777777777899888BA975BEEEAAB55689534785788888788777777755568755567667778555677788788778877777787777778877655555778777788778777765544455688875558CA655754333556655777445677655556788876885444554567555555555566677876676877654687565456775676554466776664455775456567765554557975456545455545433555565555555664434459877568757457444344345655776777777788987656788998898988888888888988888888888888888888888888888775554332333445555555443322020022223366666766777777777777777777777777777777777777777777777777899888BA975BEEEAAB55689534785788888788777777755568755567667778555677788788778877777787777778877655555778777788778777765544455688875558CA6557543335566557774456776555567888768854445545675555555555666778766768776546875654567756765544667766644557754565677655545579754565454555454335555655555556644344598775687574574443443456557767777777889876567889988989888888888889888888888888888888888888888887755543323334455555554433220200222233;
		rom_data[249] <= 3840'h7777777777777777777777777777777777777777777777778BB9898A877CEE98995478963587688887888877777855555754345567767865577777777877887677788877777777777777777778888987777887775567756887666897446865544565566677545764454456799755786556555665556656556765557875577877767775665455555555666566777654565666567654545555557B85454343324554332555555555554565555458BCA6588555578655433435555544777777888755777898899898999998989898989888898898888989888998988888765543323334445555554433222022222323666676777777777777777777777777777777777777777777777777778BB9898A877CEE98995478963587688887888877777855555754345567767865577777777877887677788877777777777777777778888987777887775567756887666897446865544565566677545764454456799755786556555665556656556765557875577877767775665455555555666566777654565666567654545555557B85454343324554332555555555554565555458BCA6588555578655433435555544777777888755777898899898999998989898989888898898888989888998988888765543323334445555554433222022222323;
		rom_data[250] <= 3840'h7777777777777777777777777777777777777777777777779A8AB98CB8AEC977877689875887987888A87777777844444432234687787777787767778877788777887777777776566777654467668998677776655666655575578AB96445665555777767777788756757766775467755765654554257764445545457765678777788867655565555667765555566567555765566543333454568855444544455543324565555555545555544479BA6555555669746633423565555887777788888A85899989989898898998988989999898899898898998989898888776544332334454555544433222202022232666767677777777777777777777777777777777777777777777777779A8AB98CB8AEC977877689875887987888A87777777844444432234687787777787767778877788777887777777776566777654467668998677776655666655575578AB96445665555777767777788756757766775467755765654554257764445545457765678777788867655565555667765555566567555765566543333454568855444544455543324565555555545555544479BA6555555669746633423565555887777788888A85899989989898898998988989999898899898898998989898888776544332334454555544433222202022232;
		rom_data[251] <= 3840'h777777777777777777777777777777777777777777777778A86BB89C88CCA8766598AA888878A77888A77777877853333234567777887777887776678777777767886677777655787775335565467788677555556754675454578877745554555557756887788777776777755556655554475566533565335544543555565667798565555667657775787755577778875566667655432334334555455577555554432367566555545555554335785454445755755543443247665466677788888997688989989989898998989989989898998989998989989988988887655443333444455554443332222022222266676677777777777777777777777777777777777777777777777778A86BB89C88CCA8766598AA888878A77888A777778778533332345677778877778877766787777777678866777776557877753355654677886775555567546754545788777455545555577568877887777767777555566555544755665335653355445435555656677985655556676577757877555777788755666676554323343345554555775555544323675665555455555543357854544457557555434432476654666777888889976889899899898989989899899898989989899989899899889888876554433334444555544433322220222222;
		rom_data[252] <= 3840'h777777777777777777777777777777777777777777777778A87CA8BB77EC8776779899788889977888877777777775454456788756756667777776777767767667777788876554567676455676555557666555656766775434677555556854455534445665677776777557766767765544557655553454345545663333577676775555666677657755677777788777675555788667544443344543455555556754432357667555555555653234553354347655555533543235776545576778797756888999999999999999989899999999899898999998998989898887665443334344545454443333222220222266666767777777777777777777777777777777777777777777777778A87CA8BB77EC87767798997888899778888777777777754544567887567566677777767777677676677777888765545676764556765555576665556567667754346775555568544555344456656777767775577667677655445576555534543455456633335776767755556666776577556777777887776755557886675444433445434555555567544323576675555555556532345533543476555555335432357765455767787977568889999999999999999898999999998998989999989989898988876654433343445454544433332222202222;
		rom_data[253] <= 3840'h7777777777777777777777777777777777777777777777779A9BA9BA69CA755799887557898A8678877777777777767776666775675555577777766776677676666678887555554555775677785443455576677756777775556765675578754565544444446767655775577788768775556565555443322454456653445886865555577765775555445555557887665544556887776555544555434454433477533333555565555655557644334334555665545445555453235557577666777975578889999999999999999999999989899999999989899899989998877655433333444444443333322222022222666676777777777777777777777777777777777777777777777777779A9BA9BA69CA755799887557898A8678877777777777767776666775675555577777766776677676666678887555554555775677785443455576677756777775556765675578754565544444446767655775577788768775556565555443322454456653445886865555577765775555445555557887665544556887776555544555434454433477533333555565555655557644334334555665545445555453235557577666777975578889999999999999999999999989899999999989899899989998877655433333444444443333322222022222;
		rom_data[254] <= 3840'h67777777777777777777777777777777777777777777777789888AB87CB87458B9797558A87875677777677877676687776676568865577777766566667767777777668765666665557555677765433345667887655557776777777756776665667555544577565444546656777577655565655554222224555555555667856645765665556555454554444345655543356557777555555454555555543334555432444455556555565576664333355567544443457834554344465775567779857777899999999999999999999999999899899999999999989998988877654433333334444343333222222222236666676667777777777777777777777777777777777777777777777789888AB87CB87458B9797558A8787567777767787767668777667656886557777776656666776777777766876566666555755567776543334566788765555777677777775677666566755554457756544454665677757765556565555422222455555555566785664576566555655545455444434565554335655777755555545455555554333455543244445555655556557666433335556754444345783455434446577556777985777789999999999999999999999999989989999999999998999898887765443333333444434333322222222223;
		rom_data[255] <= 3840'h777777777777777777777777777777777777777777777777787568A77C98645A9859857CC887557777777777776778876777777898767877677655556677666777776565565677775445544455565433444567765444566677876677677778875765567667875765433477556765554455567666542224457755555576445565577665345665675567655552335444333554356654344445555445554544543454435555555676556875555653333555654545544458544674333445655555788886557899999999999999999999999999999999998998999999999988876554333333333433333322222222222366667677777777777777777777777777777777777777777777777777787568A77C98645A9859857CC8875577777777777767788767777778987678776776555566776667777765655656777754455444555654334445677654445666778766776777788757655676678757654334775567655544555676665422244577555555764455655776653456656755676555523354443335543566543444455554455545445434544355555556765568755556533335556545455444585446743334456555557888865578999999999999999999999999999999999989989999999999888765543333333334333333222222222223;
		rom_data[256] <= 3840'h777776777777777777777777777777777777777777777778997557878B87537A6668669BA87745777778777886676A988766888888766777776555556665666766677755555545545555533444456555565555445456655556655567778889987765445568855755543576567775655577776675444356768865565444434578755565557875555556777753333444323554445442335445545445555554433456555688545796455897443455433446644467766548963565323534687455898775467899999999999999999999999999999999999999999999999998876655433333333333333233222222232366667676777776777777777777777777777777777777777777777778997557878B87537A6668669BA87745777778777886676A9887668888887667777765555566656667666777555555455455555334444565555655554454566555566555677788899877654455688557555435765677756555777766754443567688655654444345787555655578755555567777533334443235544454423354455454455555544334565556885457964558974434554334466444677665489635653235346874558987754678999999999999999999999999999999999999999999999999988766554333333333333332332222222323;
		rom_data[257] <= 3840'h667777777777777777777777777777777777777777777899CB8557868987459855888777787557777777777876778B988855677898766666777665666667676666766555455444455677777545576556545543455577667754445555677778997754455677544543556655665455555555477776555554557754455334565555787655667755556765565444544323235655545333335555544445555555434565566555556554345699655445545565445455555547A8545543453459845577875556789A999999999999999999999999999999999999999999999998877655433333333332333322222222323366666667667777777777777777777777777777777777777777777899CB8557868987459855888777787557777777777876778B988855677898766666777665666667676666766555455444455677777545576556545543455577667754445555677778997754455677544543556655665455555555477776555554557754455334565555787655667755556765565444544323235655545333335555544445555555434565566555556554345699655445545565445455555547A8545543453459845577875556789A9999999999999999999999999999999999999999999999988776554333333333323333222222223233;
		rom_data[258] <= 3840'h767677777777777777777777777777777777777777778889A9898766888755775577886567557777777777778776B987875577799877676777665567776677755677777755556556677777877655557755765556678555655555775355555788864355666634433567744788744554443446567556754355566423335566555568875434544455554444345555543566765533423356677653345445545555555445553455544333458A96555555556533454554334487554444333578645576786665689A99A9A999A999999999999999999999999999999999999999887765443332332323223233232232333366666666767677777777777777777777777777777777777777778889A9898766888755775577886567557777777777778776B987875577799877676777665567776677755677777755556556677777877655557755765556678555655555775355555788864355666634433567744788744554443446567556754355566423335566555568875434544455554444345555543566765533423356677653345445545555555445553455544333458A96555555556533454554334487554444333578645576786665689A99A9A999A9999999999999999999999999999999999999998877654433323323232232332322323333;
		rom_data[259] <= 3840'h6777677777777777777777777777777777777777778778887778985677885555675578765555787777777777877687777755677777557777767766666656676667788776655565567898665676555565556666766786554557667653444555777533575544454455555355786557776534565555556643576675333445566775578633544445555545554557755666544444322235755675432344576475665567444555555433433459B95576555578535656465333544533455346B9545575677774689AA9A999999A99A999A999999A9999999999999999999999998887655433233232232323223233233333666666676777677777777777777777777777777777777777778778887778985677885555675578765555787777777777877687777755677777557777767766666656676667788776655565567898665676555565556666766786554557667653444555777533575544454455555355786557776534565555556643576675333445566775578633544445555545554557755666544444322235755675432344576475665567444555555433433459B95576555578535656465333544533455346B9545575677774689AA9A999999A99A999A999999A9999999999999999999999998887655433233232232323223233233333;
		rom_data[260] <= 3840'h76777777777777777777777777777777777778887877788767778757669A667578678AA754578777777777778775567677777886554567776677655557657667887665456755557788986547755555555554566567888755577655532455555553345553334675544333755555667765577655444355449A75553344445657665555345445553355556765567777665333234322455334443223556664644455588545767655445544558A999A988779A888555774234444445AC545A8556676665555789AA99A9AA9A9A99A9A9A9A9999999A9A9A9A9A99999999999998877554332232232222223232323333446666666676777777777777777777777777777777777778887877788767778757669A667578678AA754578777777777778775567677777886554567776677655557657667887665456755557788986547755555555554566567888755577655532455555553345553334675544333755555667765577655444355449A75553344445657665555345445553355556765567777665333234322455334443223556664644455588545767655445544558A999A988779A888555774234444445AC545A8556676665555789AA99A9AA9A9A99A9A9A9A9999999A9A9A9A9A9999999999999887755433223223222222323232333344;
		rom_data[261] <= 3840'h77777777777777777777777777777777878877787877779888987667568879B789ACCA7554687777776778877776456567766775544566665676655556667667AA7654456655555565665556655555676544454556578765555556653345555442355555545776554445754445544434566555544333339B733324555455577654344565555554576578644458A756555434553355322222223654445544224435975555877544554454479988AA9889CCC8544554323445757CEA5597455556655444678AAA99A99A9A9A9A9A99A99A9A9A99A99A99A99A999999999998877654432222222222232323333344446666667677777777777777777777777777777777878877787877779888987667568879B789ACCA7554687777776778877776456567766775544566665676655556667667AA7654456655555565665556655555676544454556578765555556653345555442355555545776554445754445544434566555544333339B733324555455577654344565555554576578644458A756555434553355322222223654445544224435975555877544554454479988AA9889CCC8544554323445757CEA5597455556655444678AAA99A99A9A9A9A9A99A99A9A9A99A99A99A99A99999999999887765443222222222223232333334444;
		rom_data[262] <= 3840'h67767676777777777777777777777777787888788877679CBA98778756567AA78CEEB745787778777767777766675445654455555566655556655665557776779A98755556666655433455556556655766555455443467654456555553334443224555787565556556677554455534345545765553222478633335655545777754456665555565555456544459B85557545555555643343233565333443342222354543577754555445433565689888AABC85444443333456557AE87975655557654444489AA9A9A9A9AA9A9A9A99A99A9A9AA99A99A99A999999A999999887655433222222222222233333344556666666667767676777777777777777777777777787888788877679CBA98778756567AA78CEEB745787778777767777766675445654455555566655556655665557776779A98755556666655433455556556655766555455443467654456555553334443224555787565556556677554455534345545765553222478633335655545777754456665555565555456544459B85557545555555643343233565333443342222354543577754555445433565689888AABC85444443333456557AE87975655557654444489AA9A9A9A9AA9A9A9A99A99A9A9AA99A99A99A999999A99999988765543322222222222223333334455;
		rom_data[263] <= 3840'h76767676777777777777777777777788888878788777669BB9788AA7654577559EEB86778C7678766667777776565435543455555567656666655677567666777888756557777777533455558555544554556566433345554567554555322333335755776555577554566556677555566557865665223555556655544557775656657654565344343454335458875554335533456555555445443444222444333323444446556775544543357789989AAAA855544454235454348BA7657755555554455489AAAA9AA9AAAA9AA9A9A9A9A9AA9A9A9AA9AA9A9A9A999A9999887755433222222222233333334445556666667676767676777777777777777777777788888878788777669BB9788AA7654577559EEB86778C7678766667777776565435543455555567656666655677567666777888756557777777533455558555544554556566433345554567554555322333335755776555577554566556677555566557865665223555556655544557775656657654565344343454335458875554335533456555555445443444222444333323444446556775544543357789989AAAA855544454235454348BA7657755555554455489AAAA9AA9AAAA9AA9A9A9A9A9AA9A9A9AA9AA9A9A9A999A999988775543322222222223333333444555;
		rom_data[264] <= 3840'h67677777777777777777777777778778878888888777778AA89A877774357546BCA87666775687556666777775555533433556555556655776656577666666767887576567878876555555578544555444577655554334555666665555544445567755554456787653455467776457555557754565445444555543335655765556667665565433455543335445566533345653355345555444533443223434444433345435459A865444543457789899A8754455555534565333699544555555554447757AAAAAAAAAAAAAAAAAAAAA9A9A9A9AAAAAAAA99A9A99A9A99A9A988765443322222223232333344444556666667667677777777777777777777777778778878888888777778AA89A877774357546BCA87666775687556666777775555533433556555556655776656577666666767887576567878876555555578544555444577655554334555666665555544445567755554456787653455467776457555557754565445444555543335655765556667665565433455543335445566533345653355345555444533443223434444433345435459A865444543457789899A8754455555534565333699544555555554447757AAAAAAAAAAAAAAAAAAAAA9A9A9A9AAAAAAAA99A9A99A9A99A9A98876544332222222323233334444455;
		rom_data[265] <= 3840'h6667667777777777777777777878787788888887768A988AA987655554337757BB777655555576676676777765675533334755455556555777766777766666777887666757778864555654558544575555775553555433454568865655556679C9755433356777786555557644547755543455444334554457644334665555476567557766544554655544344455555555776444334434554454335443554575555755543345AC854434455445777777754434578545556433355785444455555554457679AAAAAAAAAAAAAAAAAAAAA9AAAA9AAAAAAA9A9A9A9A9A9A9A9998876544332323222232333344444555666666666667667777777777777777777878787788888887768A988AA987655554337757BB777655555576676676777765675533334755455556555777766777766666777887666757778864555654558544575555775553555433454568865655556679C9755433356777786555557644547755543455444334554457644334665555476567557766544554655544344455555555776444334434554454335443554575555755543345AC854434455445777777754434578545556433355785444455555554457679AAAAAAAAAAAAAAAAAAAAA9AAAA9AAAAAAA9A9A9A9A9A9A9A9998876544332323222232333344444555;
		rom_data[266] <= 3840'h666676767777777777777777777788888888887777AC86678755776544358777655555545557EC76677777775566553324875557777655555776787775677667787555665677775566787534544654454555455578754344456786576565567CE855653245555577555569B8555687457653343444444454433245555556556655555578776555545455544555443344457775442445333445555565455645665438A65543359A745420335644565555544434355433354543356575443345555554345668AAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAA9AAA9AAA9A9A9A9A9987655432322222232333333444455566666666666676767777777777777777777788888888887777AC86678755776544358777655555545557EC76677777775566553324875557777655555776787775677667787555665677775566787534544654454555455578754344456786576565567CE855653245555577555569B8555687457653343444444454433245555556556655555578776555545455544555443344457775442445333445555565455645665438A65543359A745420335644565555544434355433354543356575443345555554345668AAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAA9AAA9AAA9A9A9A9A99876554323222222323333334444555;
		rom_data[267] <= 3840'h777767776777777777777777788888888888887768CB76778877786457786565455433346679EB767776777656554553469754788885555567777777666667667777766676656577777765544557765655434454555455556778877755776578976665345554335554568AC96556754466533255555545553333443433456876677556798764454433455456554555445676555544444323445554554445434565368644433578656532333443453444543434433443334586347575445545555554444559AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAAA9A9A9988755433223223223333344444555566666676777767776777777777777777788888888888887768CB76778877786457786565455433346679EB767776777656554553469754788885555567777777666667667777766676656577777765544557765655434454555455556778877755776578976665345554335554568AC96556754466533255555545553333443433456876677556798764454433455456554555445676555544444323445554554445434565368644433578656532333443453444543434433443334586347575445545555554444559AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAAA9A9A99887554332232232233333444445555;
		rom_data[268] <= 3840'h67676767777777777777777877788888888888777AC978999987787557AA6775445332478777A86677667765555555555566555677765555677777676665776776678655655555776555455556655555533335443335765557777777777667777555445576553334335678997654434444544456654435444445434544555766787656677554355444545667554566545445453444555432334544444345433455445544443555545543222234333454543434543443345355237775655555555554444569BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AA9A9A98875543222222232223333445455556666666767676767777777777777777877788888888888777AC978999987787557AA6775445332478777A86677667765555555555566555677765555677777676665776776678655655555776555455556655555533335443335765557777777777667777555445576553334335678997654434444544456654435444445434544555766787656677554355444545667554566545445453444555432334544444345433455445544443555545543222234333454543434543443345355237775655555555554444569BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AA9A9A9887554322222223222333344545555;
		rom_data[269] <= 3840'h67676777777777777777777788888888888887778AB8789CCBA9778777B87776443322587777755777766765555555555544554555555556667767666666676766678765544445655443355567754444444455433355754555555555665556667555455556554222235755789753345443455557643344455555555755555565665554445453355555544455553345544332332344554542225543323345433235433444434454444454222234433455543444754574356422335875774345555665443469BAABAAAABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AA9A98876543322222222333334444555566666666767676777777777777777777788888888888887778AB8789CCBA9778777B87776443322587777755777766765555555555544554555555556667767666666676766678765544445655443355567754444444455433355754555555555665556667555455556554222235755789753345443455557643344455555555755555565665554445453355555544455553345544332332344554542225543323345433235433444434454444454222234433455543444754574356422335875774345555665443469BAABAAAABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AA9A9887654332222222233333444455556;
		rom_data[270] <= 3840'h76767677777777777777778787888888888888778A97568A99BA87779797567643422466467655677777765555548755553456534333555567766777665566677666776565555575555445555555455544467544455555444443433343455555555556755565543345564569B854555555555567544554555555555654356555545533233323454544443345532233333322222344445665335754334755544324433334344457744445422223333345432344753573458523434685575245555565455458BAAAAAAABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8876543222222222323334444455566566666676767677777777777777778787888888888888778A97568A99BA87779797567643422466467655677777765555548755553456534333555567766777665566677666776565555575555445555555455544467544455555444443433343455555555556755565543345564569B854555555555567544554555555555654356555545533233323454544443345532233333322222344445665335754334755544324433334344457744445422223333345432344753573458523434685575245555565455458BAAAAAAABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA887654322222222232333444445556;
		rom_data[271] <= 3840'h67766777777777777777778788888888888888778886656858B88875865556755564455456665677667765555555B8776556655433255555677767776555677776556656677667775676555543555554445676556555676544333223345566543454557655677545555445688755775567555575555666545544344322255555545543323224545544453233434443224443233443446765555553447865455423333333444549844435542222232333332335654433547545433475455345555555585457ABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA98875543222222222233344445555665666666767766777777777777777778788888888888888778886656858B88875865556755564455456665677667765555555B8776556655433255555677767776555677776556656677667775676555543555554445676556555676544333223345566543454557655677545555445688755775567555575555666545544344322255555545543323224545544453233434443224443233443446765555553447865455423333333444549844435542222232333332335654433547545433475455345555555585457ABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9887554322222222223334444555566;
		rom_data[272] <= 3840'h6677677777777777777777778888888888888877787789886776787655558757776676546789766666655566556678886577555553367765677776776556767775555566556775555545755555555444556766557555677643333344565455655444434543455445655455576567875444334575454567544444333233443455555555444355546655554323345544345544345444455544554454334653345443322223435556643445763223222223323454443324555444444355454356554555595447ABABAAABABABAAAAAAAAAAAAAAAAAAABABAAAAAAAAAAAAAAAAA9886553322022222223333444455556666666666677677777777777777777778888888888888877787789886776787655558757776676546789766666655566556678886577555553367765677776776556767775555566556775555545755555555444556766557555677643333344565455655444434543455445655455576567875444334575454567544444333233443455555555444355546655554323345544345544345444455544554454334653345443322223435556643445763223222223323454443324555444444355454356554555595447ABABAAABABABAAAAAAAAAAAAAAAAAAABABAAAAAAAAAAAAAAAAA9886553322022222223333444455556;
		rom_data[273] <= 3840'h6676767777777777777777888888888888888877785689777655776545577568654565557879756775555555555555664487765554566566556776666557777666553456557777555445776555655445766544555555444444434555577545554444533333333445665575566655664332344654553345434555533356555555555555455665456755544443455334576554465445543234444455333443357655333333344554334345554333334344224443334324455433554334444675555444555547ABAAABAABABABAABAAABABAAAAAABABAAAAAAAAAAAAAAAAAAAA9886543320202022233334444555556566666666676767777777777777777888888888888888877785689777655776545577568654565557879756775555555555555664487765554566566556776666557777666553456557777555445776555655445766544555555444444434555577545554444533333333445665575566655664332344654553345434555533356555555555555455665456755544443455334576554465445543234444455333443357655333333344554334345554333334344224443334324455433554334444675555444555547ABAAABAABABABAABAAABABAAAAAABABAAAAAAAAAAAAAAAAAAAA9886543320202022233334444555556;
		rom_data[274] <= 3840'h66767777777777777777777788888888888887778855775557545757987757A86655986896575567655555556545455435676545557755665566777766776566655455555555556554444555566544455543356755543333555445655565555555444433344334434445755665434433434545555432333334566454467776555665534457654465555434434333444554335753455442223323453323333467564354333444432333455433345665543233455455444544444333333556755445544455579ABBBAAAAAABAAAABBAABAAAAAAABAAAABAAAAAAAAAAAAAAAAAA8875533020202222233344455555566666666666767777777777777777777788888888888887778855775557545757987757A86655986896575567655555556545455435676545557755665566777766776566655455555555556554444555566544455543356755543333555445655565555555444433344334434445755665434433434545555432333334566454467776555665534457654465555434434333444554335753455442223323453323333467564354333444432333455433345665543233455455444544444333333556755445544455579ABBBAAAAAABAAAABBAABAAAAAAABAAAABAAAAAAAAAAAAAAAAAA887553302020222223334445555556;
		rom_data[275] <= 3840'h67677777777777777777778788888888888887777856755788545558EA669A875855877975555577555555556555543356565455468865765555677766776656765555445554444544554445555445455432347766543345775444554443455555444444545445533334445555423335544455545542222223465354335787555554434577544434433455456533433322333433233343222234443444332345453454433434222333443323355554443223465554332443355358533675555455444555579BBBBABABBBAABABAABBAABABABAAABABAAAAAAAAAAAAAAAAAAA8875533200200222333444454555566666666667677777777777777777778788888888888887777856755788545558EA669A875855877975555577555555556555543356565455468865765555677766776656765555445554444544554445555445455432347766543345775444554443455555444444545445533334445555423335544455545542222223465354335787555554434577544434433455456533433322333433233343222234443444332345453454433434222333443323355554443223465554332443355358533675555455444555579BBBBABABBBAABABAABBAABABABAAABABAAAAAAAAAAAAAAAAAAA887553320020022233344445455556;
		rom_data[276] <= 3840'h7676777777777777777788777888888888888776675787799665555AC65898755755655554755675555555556555455545544454587545666655778766777655555555545555334545775554443344533322479777544567787545555433555553444445655457875444344557543334544334334442223222344334322356454323444775345433334554457655543233454223333455433345544532334334453333444433223344333454333443334322343333223453355348533455575545445565559BBABBABABBBBABABABBAAABAAAABAAAAAABABAAAAAAAAAAAAAA987553302002022233334455555555666666767676777777777777777788777888888888888776675787799665555AC65898755755655554755675555555556555455545544454587545666655778766777655555555545555334545775554443344533322479777544567787545555433555553444445655457875444344557543334544334334442223222344334322356454323444775345433334554457655543233454223333455433345544532334334453333444433223344333454333443334322343333223453355348533455575545445565559BBABBABABBBBABABABBAAABAAAABAAAAAABABAAAAAAAAAAAAAA987553302002022233334455555555;
		rom_data[277] <= 3840'h76767777777777777777777888888888888887765679C9898555778C9668877544554543478656665555555555555665575335557754356677667887667777655555575655765454455545544333355432248B9755545677787555445546755555555545554557886554445567554434554433244333243222323344432233333333445653356533444533444655543434443333467543445444435423455543333434444542234432333554343345555422444323234664334336543345785544444455559BBBBABBBBABBBBBABBABABAABABAABAABAABAAAAAAAAAAAAAA99876543200202222334444555555556666666676767777777777777777777888888888888887765679C9898555778C9668877544554543478656665555555555555665575335557754356677667887667777655555575655765454455545544333355432248B9755545677787555445546755555555545554557886554445567554434554433244333243222323344432233333333445653356533444533444655543434443333467543445444435423455543333434444542234432333554343345555422444323234664334336543345785544444455559BBBBABBBBABBBBBABBABABAABABAABAABAABAAAAAAAAAAAAAA9987654320020222233444455555555;
		rom_data[278] <= 3840'h6777777777777777777777788888888888887775677BE9678755888B8777677545554543587556675555655555558865576455555543577778878777666677876555556655578755444444455344467533358A8555555676677775445558854565555544445545555554455556555555554444554334454233222354545322223345444433355443555443543445433434434554367433457433334324455553444544345653333332234533453537554323445333334654333334453335886544444445569BBBBBBBABBBABABABBBBABAAAABABABAAAAAAAAAAAAAAABAAAA987654322020222233444555555555666666766777777777777777777777788888888888887775677BE9678755888B8777677545554543587556675555655555558865576455555543577778878777666677876555556655578755444444455344467533358A8555555676677775445558854565555544445545555554455556555555554444554334454233222354545322223345444433355443555443543445433434434554367433457433334324455553444544345653333332234533453537554323445333334654333334453335886544444445569BBBBBBBABBBABABABBBBABAAAABABABAAAAAAAAAAAAAAABAAAA987654322020222233444555555555;
		rom_data[279] <= 3840'h7777777777777777777778888888888888887766676896468857888A875568744765565477555577565555555545875455555555434467778887877755578888755543544545776555554345555555554456665455554554556787544566654443444434458433343334455434345555433456643554443554203444445433345434443333444345765544442233233334344443343234756433244334333443444544455563322332343323554545443344535444453534332332455334886544544455558BBBBABBBBABABABBBABABBAAAABBBAAABAAABAAAABABAAAAAAA988755432020222233444555555555666666677777777777777777777778888888888888887766676896468857888A875568744765565477555577565555555545875455555555434467778887877755578888755543544545776555554345555555554456665455554554556787544566654443444434458433343334455434345555433456643554443554203444445433345434443333444345765544442233233334344443343234756433244334333443444544455563322332343323554545443344535444453534332332455334886544544455558BBBBABBBBABABABBBABABBAAAABBBAAABAAABAAAABABAAAAAAA988755432020222233444555555555;
		rom_data[280] <= 3840'h666777777777777777778888888888888888777566565555755A879986557975665588555555666656555555555875555445545544567788877787765557889886544332455444554555434544555443457753333334544344455555445445433333334458B523222234456423344554334445434554433554224433345554455334543234433456775434433222234455444332222225655443333333322233334444564464443333553225653443333433456444453354323334355434675644544455557ABABBABBBBBAABAABBABABBBABAABBBAAABABABAAABABAAAAAAA9877553322222233344555555555566666666666777777777777777778888888888888888777566565555755A879986557975665588555555666656555555555875555445545544567788877787765557889886544332455444554555434544555443457753333334544344455555445445433333334458B523222234456423344554334445434554433554224433345554455334543234433456775434433222234455444332222225655443333333322233334444564464443333553225653443333433456444453354323334355434675644544455557ABABBABBBBBAABAABBABABBBABAABBBAAABABABAAABABAAAAAAA98775533222222333445555555555;
		rom_data[281] <= 3840'h7777777777777777777878888888888888887766755557A7558A76898545996575558755543555555555555545559544554556457875778778888755555778A8755543234775333344533444444433334565434433354333433332344433334444444455568532332344467545554555455433335654445643344443456654443356644443344555554444444322235786555533432333333333334433432322334544543555654333443335534433334333356323333365323337534553455544444445557ABBBBBBBABBBBBBBABAAABBAABBBABABABABBABAAAAAABAAAAAA98876553322222233444555555555666666667777777777777777777878888888888888887766755557A7558A76898545996575558755543555555555555545559544554556457875778778888755555778A8755543234775333344533444444433334565434433354333433332344433334444444455568532332344467545554555455433335654445643344443456654443356644443344555554444444322235786555533432333333333334433432322334544543555654333443335534433334333356323333365323337534553455544444445557ABBBBBBBABBBBBBBABAAABBAABBBABABABABBABAAAAAABAAAAAA98876553322222233444555555555;
		rom_data[282] <= 3840'h67676767777777777777878888888888888887657577689857A8557996569844556777655345555555555545555485455566775566557887788887655577777755455335444334444443455444444334445544455543223333332334345433433344545554554345455545775675555555454334443334543356445544554345544554453344333334434456442233456556753333334322222234543244322345764233454454323323323434444435535534556523433233334A534643555544443455557ABABABBBBBBBBBBBBBBBABABAAABBBABBBAABBAAABABAAAABAAA988876553322223334455555555556666667667676767777777777777878888888888888887657577689857A8557996569844556777655345555555555545555485455566775566557887788887655577777755455335444334444443455444444334445544455543223333332334345433433344545554554345455545775675555555454334443334543356445544554345544554453344333334434456442233456556753333334322222234543244322345764233454454323323323434444435535534556523433233334A534643555544443455557ABABABBBBBBBBBBBBBBBABABAAABBBABBBAABBAAABABAAAABAAA98887655332222333445555555555;
		rom_data[283] <= 3840'h66776777777777777787888888888888888887767687567769854468A55786434665677555565555565555555543544555577657865677667778875556787777555454575334444543345554457765433334554455543333332334454575555435555433443554555555445776555455544554444333432223455553355544555433323345533322333434443343443233344433433553222202554335333223446533355444534433243323334435543354333333233433233468334544455543554455458ABABBBBBBBBBBABBBBBBBBBBBBBBBBBBABBBABABAAAAABAAAAAAA99887654432232334555555666666667666766776777777777777787888888888888888887767687567769854468A55786434665677555565555565555555543544555577657865677667778875556787777555454575334444543345554457765433334554455543333332334454575555435555433443554555555445776555455544554444333432223455553355544555433323345533322333434443343443233344433433553222202554335333223446533355444534433243323334435543354333333233433233468334544455543554455458ABABBBBBBBBBBABBBBBBBBBBBBBBBBBBABBBABABAAAAABAAAAAAA9988765443223233455555566666;
		rom_data[284] <= 3840'h77677777777777777778888888888888888887667577556667643468944545555875576555545555565555554556445775445537875656667777887555777766555434455443434334565454479985445555433444434443233444454454577545654454443333345565444664445445444675444444432333234432575444443332223355444543233443333343334322223223333433332232453355322343334333455433345432344544434345432343434433543343333555354457446443563455457ABBBBBBBBBBBBBBABABABBBBBBBBABABABABBBBAAAABAABAAAABAA9987765433323344555555565666666667677677777777777777778888888888888888887667577556667643468944545555875576555545555565555554556445775445537875656667777887555777766555434455443434334565454479985445555433444434443233444454454577545654454443333345565444664445445444675444444432333234432575444443332223355444543233443333343334322223223333433332232453355322343334333455433345432344544434345432343434433543343333555354457446443563455457ABBBBBBBBBBBBBBABABABBBBBBBBABABABABBBBAAAABAABAAAABAA998776543332334455555556566;
		rom_data[285] <= 3840'h667767777777777777887888888888888888877775787556575323688433344478745667755555555655555555574347753443567655556666677755556777655554334344434554345753334777654565555444332355433233333434345554444333454333333434545445433355654557754343433233332222025543444433443354334434433344443335554333322222232332202323323434754433333333445544543343344445432354333333323234334433432223454554554454335634565579BBABBBBBBBBABBBABABBABABABABBBBBBBBBBABABAAAAAAAAAAAAAA987665443233444555566666666676666667767777777777777887888888888888888877775787556575323688433344478745667755555555655555555574347753443567655556666677755556777655554334344434554345753334777654565555444332355433233333434345554444333454333333434545445433355654557754343433233332222025543444433443354334434433344443335554333322222232332202323323434754433333333445544543343344445432354333333323234334433432223454554554454335634565579BBABBBBBBBBABBBABABBABABABABBBBBBBBBBABABAAAAAAAAAAAAAA9876654432334445555666666;
		rom_data[286] <= 3840'h777777777777777778778888888888888888877775687655567334776335555576644665555555555555555555564445545333567765577666777555556776544344444345444544334443233445444453455443322467543332344433444333332333355444554555455544433444534566543343333333342000233333455543443333223543333565454434765433333022554333322334433333544553354434446754444233344333233454332223322333343333332232344674345544435534567669BBABBBBBBBBBBBBBBBBBBBABABBABBABAABABBABAAAABABAAAAAAAAA88775543333445555666666666667677777777777777777778778888888888888888877775687655567334776335555576644665555555555555555555564445545333567765577666777555556776544344444345444544334443233445444453455443322467543332344433444333332333355444554555455544433444534566543343333333342000233333455543443333223543333565454434765433333022554333322334433333544553354434446754444233344333233454332223322333343333332232344674345544435534567669BBABBBBBBBBBBBBBBBBBBBABABBABBABAABABBABAAAABABAAAAAAAAA887755433334455556666666;
		rom_data[287] <= 3840'h767677777777777787878888888888889888887765565675567335654225555557734544456555555645555545555644335433457665677656777555557665443334443457653333543233333244445533334343333567543433455434554333333454445556754575576555433444343344323344333334333222232345454543334444333443234664343332454333443223675435533346443322233333454445335543233223333322333353343344233333333443343233343553357555434433456558BBBBBBBBBBBBBBBBBBBABABABBBBBBBABBBBBAAAAAAAAAAAAABAAAAA98877654433445555666666666676767767677777777777787878888888888889888887765565675567335654225555557734544456555555645555545555644335433457665677656777555557665443334443457653333543233333244445533334343333567543433455434554333333454445556754575576555433444343344323344333334333222232345454543334444333443234664343332454333443223675435533346443322233333454445335543233223333322333353343344233333333443343233343553357555434433456558BBBBBBBBBBBBBBBBBBBABABABBBBBBBABBBBBAAAAAAAAAAAAABAAAAA988776544334455556666666;
		rom_data[288] <= 3840'h676777777777777777787888888888888888887765777875574335543234345446544445456545555555555555456863334445556665678655667765556555545444344356653334653223553245445535432333343444434544453234444554344466435667544555587567544544554223233444344444334323333355454532344567553333433333333432223234433334444334332345433332222223233344234432223323223323334333355543345333333563254345644433456555444433356559CBBBBBBBBBBBBBBBBABBBBAAABABABABABBABBBAAABABABABAAAAAAAAA887655444445555667776666666666676777777777777777787888888888888888887765777875574335543234345446544445456545555555555555456863334445556665678655667765556555545444344356653334653223553245445535432333343444434544453234444554344466435667544555587567544544554223233444344444334323333355454532344567553333433333333432223234433334444334332345433332222223233344234432223323223323334333355543345333333563254345644433456555444433356559CBBBBBBBBBBBBBBBBABBBBAAABABABABABBABBBAAABABABABAAAAAAAAA8876554444455556677766;
		rom_data[289] <= 3840'h676767777777777787888888888888888988887777878977753344553364345433445555555445555556754555545765335555555655577655557776555555555543456544444444443335665335443445544443333333223333433232333444333456433455433455575556555444664222335554345653345334544444344333344455544433433222334553202224334433222222223433422333320222323243235543224333443334344333234432355433332343344346974435534554444333457569BBBBBBBBBBBBBABBBBBBBBBBBABBBBABBBABBABBBBAAABAABABAAAAAA9987765544445555666767766676666676767777777777787888888888888888988887777878977753344553364345433445555555445555556754555545765335555555655577655557776555555555543456544444444443335665335443445544443333333223333433232333444333456433455433455575556555444664222335554345653345334544444344333344455544433433222334553202224334433222222223433422333320222323243235543224333443334344333234432355433332343344346974435534554444333457569BBBBBBBBBBBBBABBBBBBBBBBBABBBBABBBABBABBBBAAABAABABAAAAAA99877655444455556667677;
		rom_data[290] <= 3840'h767677777777777777888888888888888989887778777757745445555564489444656543343445555555555555444554446653665566665655555655555544454343455543333544334346565434433333455554332222333433443333333433343445422333223554454445555444444333434553323443333233543333343333334423333434433323333544200232256433222232235302222333332233343332245433224333465533333443322323443343333233332336A85335534554434333455569BBBBBBBBBBBABBBBBBBBBABBBBBABBBABBBABBBABABBABBAAAAAAABABA998775555445555566667666667667767677777777777777888888888888888989887778777757745445555564489444656543343445555555555555444554446653665566665655555655555544454343455543333544334346565434433333455554332222333433443333333433343445422333223554454445555444444333434553323443333233543333343333334423333434433323333544200232256433222232235302222333332233343332245433224333465533333443322323443343333233332336A85335534554434333455569BBBBBBBBBBBABBBBBBBBBABBBBBABBBABBBABBBABABBABBAAAAAAABABA9987755554455555666676;
		rom_data[291] <= 3840'h666676777777777788888888888888988998877777666544545468678333698554535532333456555555555444543345545775665677665666644445565544323333433324443444433355343333334322334565644433355554335543456643355555532222233444433344444443323454322332220202202232333223554333335642222233235533333222332223455334533233333022222224745334542332223233222222344322432343222233322453243233332455633444334545443333445559CBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBABBBBBABABAAAABABAABAA98876555445555555667666666676666676777777777788888888888888988998877777666544545468678333698554535532333456555555555444543345545775665677665666644445565544323333433324443444433355343333334322334565644433355554335543456643355555532222233444433344444443323454322332220202202232333223554333335642222233235533333222332223455334533233333022222224745334542332223233222222344322432343222233322453243233332455633444334545443333445559CBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBABBBBBABABAAAABABAABAA988765554455555556676;
		rom_data[292] <= 3840'h677767777777777778788888888888989898877776797544435556555433688655754344443555555555555445454456875554445776565556544455555444323333323235543434443344432344333223443334444333234554454345567743377644333222234455344555544343223564333223332002232333222234553454345753322443347653332222333323322235322332232020202235533345432323553233332233323234333344433232323354344332325633544323333455444343445558BBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBABABABABBBBABBBABAABAABA99877655444445555556666666767677767777777777778788888888888989898877776797544435556555433688655754344443555555555555445454456875554445776565556544455555444323333323235543434443344432344333223443334444333234554454345567743377644333222234455344555544343223564333223332002232333222234553454345753322443347653332222333323322235322332232020202235533345432323553233332233323234333344433232323354344332325633544323333455444343445558BBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBABABABABBBBABBBABAABAABA998776554444455555566;
		rom_data[293] <= 3840'h6666777777777778888888888888898989988878759C9676545875443555567545744456674445454555554444434558C85554344655655555554555555444334433343344333555544333323345544343433322232334322334543345555543455543343332344454544544444443335543333223433332333433220354333454444433344543335754233223333333222233223333320222002333322233323333543333332233223333355333533223345333234322324533455333343344443343355458CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABABAABAAABBA98776555444444455555666676666666777777777778888888888888898989988878759C9676545875443555567545744456674445454555554444434558C85554344655655555554555555444334433343344333555544333323345544343433322232334322334543345555543455543343332344454544544444443335543333223433332333433220354333454444433344543335754233223333333222233223333320222002333322233323333543333332233223333355333533223345333234322324533455333343344443343355458CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABABAABAAABBA98776555444444455555;
		rom_data[294] <= 3840'h6666667777777777788888888888888899898878759A7688654774433655456535633455453444545555444443345656875444345677555554555455555545444434555432234555433322334555443454333443223345533223433334434332334332356653334444444445544334333233344233333333223323222354233554443455446543334553344333223333322320234323222223223322202322234333333233222222222345456533432443343233233353323333354334444353443443345558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBABBABABABBBABBAAAAAABABAAAA9877554434334344455666666676666667777777777788888888888888899898878759A7688654774433655456535633455453444545555444443345656875444345677555554555455555545444434555432234555433322334555443454333443223345533223433334434332334332356653334444444445544334333233344233333333223323222354233554443455446543334553344333223333322320234323222223223322202322234333333233222222222345456533432443343233233353323333354334444353443443345558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBABBABABABBBABBAAAAAABABAAAA9877554434334344455;
		rom_data[295] <= 3840'h666676777777777787888888888898989898888877987667554786554534345434535554342444554554544434555655765554655676555554555455554568655443455432233443333323335543343455334554335433333222334333332333233322457744334333455657743345432234333333333422343234323432333354344443334533444443334332233233223322234322233333334322222320355333323222222232233345555533232443232343333344424423344434434354433443444568CBBBBBBBBBBBABBBBBBBBBBBBBBABBBBBBBBABBBBBBABBBAAAABABBAAABAA988765433333333344566666676666676777777777787888888888898989898888877987667554786554534345434535554342444554554544434555655765554655676555554555455554568655443455432233443333323335543343455334554335433333222334333332333233322457744334333455657743345432234333333333422343234323432333354344443334533444443334332233233223322234322233333334322222320355333323222222232233345555533232443232343333344424423344434434354433443444568CBBBBBBBBBBBABBBBBBBBBBBBBBABBBBBBBBABBBBBBABBBAAAABABBAAABAA9887654333333333445;
		rom_data[296] <= 3840'h76666676777777777888888888888989999988888987774455477776445434535543654433244545454454443455344576555565556575545554455555457A755433333333322333455333233333332333334433345432322222224543444433332223455434434433567888533354434443232334553333344334334433343234333233432223332322222332233433334433232222343322323333332223554233334323234443334333434433232342223333233223344422344444344444443333345558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBABBBAAABBBBABA98876543322322333446666766676666676777777777888888888888989999988888987774455477776445434535543654433244545454454443455344576555565556575545554455555457A755433333333322333455333233333332333334433345432322222224543444433332223455434434433567888533354434443232334553333344334334433343234333233432223332322222332233433334433232222343322323333332223554233334323234443334333434433232342223333233223344422344444344444443333345558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBABBBAAABBBBABA9887654332232233344;
		rom_data[297] <= 3840'h667677777777777787888888888889899898888889777555555445653475455597445444534344445545544444333233445543444555655555554445555457755532322243333234454443222334433322233222233333332322223664476433333333333237545653455775323343343442333457752223223333234444453223222245432343222220222223234544565543332222345220203444322225533334333235445544544323333333233332323223232324244323343443335434433333446558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBABABBBABABABABAABA988755432222222333466666666667677777777777787888888888889899898888889777555555445653475455597445444534344445545544444333233445543444555655555554445555457755532322243333234454443222334433322233222233333332322223664476433333333333237545653455775323343343442333457752223223333234444453223222245432343222220222223234544565543332222345220203444322225533334333235445544544323333333233332323223232324244323343443335434433333446558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBABABBBABABABABAABA9887554322222223334;
		rom_data[298] <= 3840'h666767777777777778888888888889989989888877576576675434443454333795654345545444555544444443333334434434434554555545555445555545555444433234443344332354232355542223333233223333233333224554344333333333332346557754334543233333333233335677633224334753335444463222222465433553222020232223323234754332334223255322235432232233322323222255333323553422333233323333322233334433333433433433234535443333346559CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBBABBBAAABAA988755333222222223366666666666767777777777778888888888889989989888877576576675434443454333795654345545444555544444443333334434434434554555545555445555545555444433234443344332354232355542223333233223333233333224554344333333333332346557754334543233333333233335677633224334753335444463222222465433553222020232223323234754332334223255322235432232233322323222255333323553422333233323333322233334433333433433433234535443333346559CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBBABBBAAABAA9887553332222222233;
		rom_data[299] <= 3840'h666767677777777788888888888898999898888777676565454443433433323786543343445344555544444443355345544567445554558755554444555545555445543334554333333433333343332225532343333333234532232333343245522332222334455554333332234555333222333433333234445885445544763222222454333543323222332223322223432202233222244232345322233322223222322254222223433533343332334323332333334542233344433443333435543333445558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBABBBABBBBABA998755332222222223366666666666767677777777788888888888898999898888777676565454443433433323786543343445344555544444443355345544567445554558755554444555545555445543334554333333433333343332225532343333333234532232333343245522332222334455554333332234555333222333433333234445885445544763222222454333543323222332223322223432202233222244232345322233322223222322254222223433533343332334323332333334542233344433443333435543333445558CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBABBBABBBBABA9987553322222222233;
		rom_data[300] <= 3840'h66666677777777777888888888989898999888877765556445465553333544457774454574554555554444544336855754455533455456775565444457745544343443222345533334455333332222233443334343355542355333223343335543223222333433343323233333567653232333222202333332355544333454322222323223333334432223223322232232022222002344423223443232222223223332223322223433553244433486334423344433324233333444444345443554333335655ACBBBBCBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBAA99876542322222222236666666666666677777777777888888888989898999888877765556445465553333544457774454574554555554444544336855754455533455456775565444457745544343443222345533334455333332222233443334343355542355333223343335543223222333433343323233333567653232333222202333332355544333454322222323223333334432223223322232232022222002344423223443232222223223332223322223433553244433486334423344433324233333444444345443554333335655ACBBBBCBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBAA9987654232222222223;
		rom_data[301] <= 3840'h66677776777777777788888888889898988988886886566443575455335644576664542343444454555444544344544565435322445455555555444457645554333232333334443443367544222222232334432222345542356554322454344432223323554333332222222333335542322222332000020002343443222223233222322234430477534333255323443222033222222343323223432233000233442233222234442333433345423576444333233234323223333343443444344443334345745ABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABABBBABABBABAA8876543232222222326666666666677776777777777788888888889898988988886886566443575455335644576664542343444454555444544344544565435322445455555555444457645554333232333334443443367544222222232334432222345542356554322454344432223323554333332222222333335542322222332000020002343443222223233222322234430477534333255323443222033222222343323223432233000233442233222234442333433345423576444333233234323223333343443444344443334345745ABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABABBBABABBABAA887654323222222232;
		rom_data[302] <= 3840'h666676777777777778888888888899989898888779855556565466575455555764545764533544444555544443443344544444334455555544544444555455444433323333332333333555332323323232234322222243233577642223332323223232355542222233542223432233222234233344433220023322224433223432333323343335543345334543235533333222232222222222243322322222233323433222234422355333344335754443322323443233232354353334344555543333455459CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBBABBABBBBABAAAA88755432323222223266666666666676777777777778888888888899989898888779855556565466575455555764545764533544444555544443443344544444334455555544544444555455444433323333332333333555332323323232234322222243233577642223332323223232355542222233542223432233222234233344433220023322224433223432333323343335543345334543235533333222232222222222243322322222233323433222234422355333344335754443322323443233232354353334344555543333455459CBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBBABBABBBBABAAAA887554323232222232;
		rom_data[303] <= 3840'h66666777777778788888888888989899898888877854555788546755555455675554585463564344555454443344444433343544344555554455545444554455554433344322233333344333333233234334443323333223445643223343333232223344442233333344323343222002332222355785432222333333443322333444543343333322023333333224543333222222243200000234432333223322322542223322332347534323322453334322232343323333225534434444555754333344446ACBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBABBABBBBABAA9876543232322222236666666666666777777778788888888888989899898888877854555788546755555455675554585463564344555454443344444433343544344555554455545444554455554433344322233333344333333233234334443323333223445643223343333232223344442233333344323343222002332222355785432222333333443322333444543343333322023333333224543333222222243200000234432333223322322542223322332347534323322453334322232343323333225534434444555754333344446ACBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBABBABBBBABAA987654323232222223;
		rom_data[304] <= 3840'h66666667777777787888888888888989898888876654555566545644455435555555553353675334455444554345454323444554444545544454544434554565554433343333323553233344344223233323443332332223333322222344554222323333222233433333333433222223443222345564333222333432233333334665543343332002222342222233332322223422244322220224432343222223223432235422222346443322223532334322233233332232024444344445554554343334446ACBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBABBBAA99876543323232322226666666666666667777777787888888888888989898888876654555566545644455435555555553353675334455444554345454323444554444545544454544434554565554433343333323553233344344223233323443332332223333322222344554222323333222233433333333433222223443222345564333222333432233333334665543343332002222342222233332322223422244322220224432343222223223432235422222346443322223532334322233233332232024444344445554554343334446ACBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBABBBAA9987654332323232222;
		rom_data[305] <= 3840'h66667677777777778788888888899989988888875665455556534663344344445476323454564344454444454345433333455454444455445545534345544554443233233343334433332333344233422223332332222222223222222234543223432222222323443343333334432222354332322322022333322322245454335775543233433333233443332332333322225532233222222223322453322222334320224322222344443220234443333323322322323232222334344345444443333344546ACBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBBBABABBBBAAAAA9886543323222222235556666666667677777777778788888888899989988888875665455556534663344344445476323454564344454444454345433333455454444455445545534345544554443233233343334433332333344233422223332332222222223222222234543223432222222323443343333334432222354332322322022333322322245454335775543233433333233443332332333322225532233222222223322453322222334320224322222344443220234443333323322322323232222334344345444443333344546ACBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBBBABABBBBAAAAA988654332322222223;
		rom_data[306] <= 3840'h66666677777777878888888889888998988888876785478857534884432344544375323554354433444544454445433444355533555455545555534355434343233223333232245322333222233345532222222353202332222022433223332333443222222232345443543334443232222223222000202322202023346775434553332344323544332323554433233322334322300002232333323443432223332222232222023343443222223333333345222333223224332035433335554443333344447BCCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBABA9987554332222222226565656666666677777777878888888889888998988888876785478857534884432344544375323554354433444544454445433444355533555455545555534355434343233223333232245322333222233345532222222353202332222022433223332333443222222232345443543334443232222223222000202322202023346775434553332344323544332323554433233322334322300002232333323443432223332222232222023343443222223333333345222333223224332035433335554443333344447BCCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBABA998755433222222222;
		rom_data[307] <= 3840'h66666767777777788888888888999898988888876787578555425975433436853454554344544444344444434343455555334324565555555455433444455543333333323223244322332343332333332203333223223443222234433223232233433245423322223334653232222332020022220202222220022223323553243333323344233332222333455332323323322022200023432333322222220244222322332222223232232322322343333322323333223232332235444334555443333445437CCBBBBBBBBBCBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBBBBBBABABA9977553322222222235656666666666767777777788888888888999898988888876787578555425975433436853454554344544444344444434343455555334324565555555455433444455543333333323223244322332343332333332203333223223443222234433223232233433245423322223334653232222332020022220202222220022223323553243333323344233332222333455332323323322022200023432333322222220244222322332222223232232322322343333322323333223232332235444334555443333445437CCBBBBBBBBBCBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBBBBBBABABA997755332222222223;
		rom_data[308] <= 3840'h66666677777777778888888888889899888888875755776555348854546535743653565445543455545444443445654333334235885544567555434333455443333234335322333333322343234332223233332222232333333232222334443333332357543322222034443222222202232223332233223222232223332223233333323323332223322332233223333333432202022222224323222002002355222220222322223322233222202323334423333333222222443324344334554443333444447BCBBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBABBBAAAA877553322222022225656666666666677777777778888888888889899888888875755776555348854546535743653565445543455545444443445654333334235885544567555434333455443333234335322333333322343234332223233332222232333333232222334443333332357543322222034443222222202232223332233223222232223332223233333323323332223322332233223333333432202022222224323222002002355222220222322223322233222202323334423333333222222443324344334554443333444447BCBBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBABBBAAAA87755332222202222;
		rom_data[309] <= 3840'h66676777777777788888888889999998888888776554555556578755546546755644544554433355545344454444444433453347765554567754344334455443432233334323232345334323454320222332220023333223333322224435554332322344433322222222322222232332223244432222224322233325532202232233334334543344223322222002233322222220234202003222220202022333223220222222223332223222022223343333344323222220233334334334445444333444448CCBBBBBBBBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABABA9887543222222222225566566666676777777777788888888889999998888888776554555556578755546546755644544554433355545344454444444433453347765554567754344334455443432233334323232345334323454320222332220023333223333322224435554332322344433322222222322222232332223244432222224322233325532202232233334334543344223322222002233322222220234202003222220202022333223220222222223332223222022223343333344323222220233334334334445444333444448CCBBBBBBBBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABABA988754322222222222;
		rom_data[310] <= 3840'h6667667777777878888888889889998988888878665556544468767654455444555555458333334554434555444543344433336A965654454444455533344443454333433343323343344323333322233320223222233323334322223334433322222233323332322222222022232333222233322022222232344235422003332355543334322443233332020023333232200020223202322023202202202222355222222222222222022223222422343323333333332233332343233334445443344354458CBCBBCBBBBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBABBAAA88754322020020222655665666667667777777878888888889889998988888878665556544468767654455444555555458333334554434555444543344433336A965654454444455533344443454333433343323343344323333322233320223222233323334322223334433322222233323332322222222022232333222233322022222232344235422003332355543334322443233332020023333232200020223202322023202202202222355222222222222222022223222422343323333333332233332343233334445443344354458CBCBBCBBBBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBABBAAA88754322020020222;
		rom_data[311] <= 3840'h6666677777777788788888888999999889888888666567753355677543454543434455346453333555434445544553235643446B955554444333469754434432334333432444232232233323222222345322224432222244323322222223222202022222322454222343222320222344432223333233320202233233222233222346543322235433234422200233332232002222202023320024220020002332365344202220200022222233332332433332222222322343322342344443465554333444458CBBBBBCBCBCBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABABABBABA998754332202202222565656666666677777777788788888888999999889888888666567753355677543454543434455346453333555434445544553235643446B955554444333469754434432334333432444232232233323222222345322224432222244323322222223222202022222322454222343222320222344432223333233320202233233222233222346543322235433234422200233332232002222202023320024220020002332365344202220200022222233332332433332222222322343322342344443465554333444458CBBBBBCBCBCBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABABABBABA998754332202202222;
		rom_data[312] <= 3840'h66676777777777788888888898989999888888886555567544445764324445544233553355644334544444445434334345544458754444444434467554333432222233333344323223222233220223343322333342222244332232222222222022202002223685322355345532002234332023443223222200222322223442222223332322245333344322222232222223222223320222220233223332203532354453222222222200233333222233333233222222222333323333334443457543433443359CCCCCBCBCBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABA9987553222200222236556666666676777777777788888888898989999888888886555567544445764324445544233553355644334544444445434334345544458754444444434467554333432222233333344323223222233220223343322333342222244332232222222222022202002223685322355345532002234332023443223222200222322223442222223332322245333344322222232222223222223320222220233223332203532354453222222222200233333222233333233222222222333323333334443457543433443359CCCCCBCBCBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABA998755322220022223;
		rom_data[313] <= 3840'h66766777777777888888888899999999888888886534444545535565234344555443554355433333444444344333334443334334555445544444354333444443222333222233334322222233222222233233320222333323333232222334432222222022223685322246677653220222222222233222023202203323433332223222022333322223345422223332223223222003320223222233333442023433443432222332322202432232222223322233323333222322333232233344457533333444359CCBBCBBCBCBBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABAAABA9987543320222022225566656666766777777777888888888899999999888888886534444545535565234344555443554355433333444444344333334443334334555445544444354333444443222333222233334322222233222222233233320222333323333232222334432222222022223685322246677653220222222222233222023202203323433332223222022333322223345422223332223223222003320223222233333442023433443432222332322202432232222223322233323333222322333232233344457533333444359CCBBCBBCBCBBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABAAABA998754332022202222;
		rom_data[314] <= 3840'h6666677777778787888888888989999988888888764344543544566535433344555354324532333334343443333334444233233334444655444443434345545532333333220223332222233332222223223322222223222244323222334555222333222222234320222456554322202020223222322222222222232354223233333020233222232224753222332232322222020220023332223232232222223333322222333332222233232322222232322333332222223223333233333445654333344536ACCCCBCCBCBCCBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBABAA98765322020022223556566666666677777778787888888888989999988888888764344543544566535433344555354324532333334343443333334444233233334444655444443434345545532333333220223332222233332222223223322222223222244323222334555222333222222234320222456554322202020223222322222222222232354223233333020233222232224753222332232322222020220023332223232232222223333322222333332222233232322222232322333332222223223333233333445654333344536ACCCCBCCBCBCCBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBABAA98765322020022223;
		rom_data[315] <= 3840'h6666677777777788888888989899999888888888764434533434467535333343334333334542234333333443333333433342345433345555444434343343455433333234320202322233335533332333222332222233322335322322344343222345322022222232022233332220002022245433422000002222222333223232232202233323442223554320202222222320002000002220223222222220022222222234333333333432323322322332332223333222233222333233454345554333344447BCCBCBCBCBCBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBAA98765432202202223555665666666677777777788888888989899999888888888764434533434467535333343334333334542234333333443333333433342345433345555444434343343455433333234320202322233335533332333222332222233322335322322344343222345322022222232022233332220002022245433422000002222222333223232232202233323442223554320202222222320002000002220223222222220022222222234333333333432323322322332332223333222233222333233454345554333344447BCCBCBCBCBCBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBAA98765432202202223;
		rom_data[316] <= 3840'h6667667777777778888888889899998988888888754444533433457523343235433334334543333333333343333233323433355333445554443344344434465333333333223322222353334323323542222234323544322343222323432220202333202220222443222222222002200223357533320000002333332222343332322232245422332223344443224522332320022000200000023200223332222222220233333233333233323333333233442002333223332223322223433454444333344347BCCBCBCBCBCBCBBCCCCBCCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABBA99875432220022222656566666667667777777778888888889899998988888888754444533433457523343235433334334543333333333343333233323433355333445554443344344434465333333333223322222353334323323542222234323544322343222323432220202333202220222443222222222002200223357533320000002333332222343332322232245422332223344443224522332320022000200000023200223332222222220233333233333233323333333233442002333223332223322223433454444333344347BCCBCBCBCBCBCBBCCCCBCCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABBA99875432220022222;
		rom_data[317] <= 3840'h6666777777777878888888898999999888888888775455534554456434433334434344333553333333333344333355333333343323444554443443334333344334422222222222223430222322222322332334323653222222222222222222202202223222345532302222222003322232333322220023222223332222323323222222243223322222223443233222320222220000202022233320234222222023322233323223332332344222234432332223222223233223322444443453333333444448BCBCBCBCBCBCBCCBBBBCBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABAA9876432202202223555666666666777777777878888888898999999888888888775455534554456434433334434344333553333333333344333355333333343323444554443443334333344334422222222222223430222322222322332334323653222222222222222222202202223222345532302222222003322232333322220023222223332222323323222222243223322222223443233222320222220000202022233320234222222023322233323223332332344222234432332223222223233223322444443453333333444448BCBCBCBCBCBCBCCBBBBCBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABAA9876432202202223;
		rom_data[318] <= 3840'h6667667777777888888888898989999888888888755555554555434243344664335344322464333233323343333356433454332334334443343443343333334333322323342202245322022220202222453233433432223220200202202020220222332223433222220222222022332222022222222233332220202332334223322332222223222234422222222222202320233202322020333022333222222223322322323222332233443222224653232223202202233233223534333445433333443448CCCBCBCBCBCBCBBCCCCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA99876543200202222555555666667667777777888888888898989999888888888755555554555434243344664335344322464333233323343333356433454332334334443343443343333334333322323342202245322022220202222453233433432223220200202202020220222332223433222220222222022332222022222222233332220202332334223322332222223222234422222222222202320233202322020333022333222222223322322323222332233443222224653232223202202233233223534333445433333443448CCCBCBCBCBCBCBBCCCCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA99876543200202222;
		rom_data[319] <= 3840'h6666676777777788888888898999999888888887755455674544332243355555534278534354332333232333333334333575322343244454334433343333343433233433442222243332233332000222343222222222222222202222022022202234532022222022220202022002222022222222233232202200233233323222233232222232202255322202020222223220222334320202222222333222233323333223223222222333543333223654323222022222222343223333433335433333434359CBCCCCBCBCBCBCCBBBBBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABABAA9887543220022223555566666666676777777788888888898999999888888887755455674544332243355555534278534354332333232333333334333575322343244454334433343333343433233433442222243332233332000222343222222222222222202222022022202234532022222022220202022002222022222222233232202200233233323222233232222232202255322202020222223220222334320202222222333222233323333223223222222333543333223654323222022222222343223333433335433333434359CBCCCCBCBCBCBCCBBBBBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABABAA9887543220022223;
		rom_data[320] <= 3840'h66676777777777888888888989999999888888877545557645555334333533344443AB546443323333233233233333323554333333245554334444333334433433344332322202222322244322020202220000202234322222222222223222234555432202202220223302243220202003454323332222222022222222222222232023432322002343332222232233332222220233220020022322223223244323232022233232232233443433223543333223222222222343223333433434433443344349CCCBCBCCCCCCCBBCCCCCBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABA9875532220002225565556666676777777777888888888989999999888888877545557645555334333533344443AB546443323333233233233333323554333333245554334444333334433433344332322202222322244322020202220000202234322222222222223222234555432202202220223302243220202003454323332222222022222222222222232023432322002343332222232233332222220233220020022322223223244323232022233232232233443433223543333223222222222343223333433434433443344349CCCBCBCCCCCCCBBCCCCCBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABA987553222000222;
		rom_data[321] <= 3840'h666676777777778888888888999999988888888775455555466455443443322333348954443322332232333233333332354333333234554333344333334344333334422222220222322223322220202222222222444542223222022222222023443332203322334324553245532002022345222355300022022202232332233222022333332235232233322223223222202342000000000022332223223223222233222223233223222333432222334333222232222222323322333334434443343344435ACCBCBCBCBBCBBCCBBBBBBBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBA99765432002222255555556666676777777778888888888999999988888888775455555466455443443322333348954443322332232333233333332354333333234554333344333334344333334422222220222322223322220202222222222444542223222022222222023443332203322334324553245532002022345222355300022022202232332233222022333332235232233322223223222202342000000000022332223223223222233222223233223222333432222334333222232222222323322333334434443343344435ACCBCBCBCBBCBBCCBBBBBBBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBA997654320022222;
		rom_data[322] <= 3840'h666667777777787888888888889999998888788875556555355355323344433233235663223333222332232222333333233322223333543333344333333334434432232222202243222023223222022222223323333222223222223220202022222220002222344334433345532222222222222355322200222300332333333220033223433555322223322320220222220330000000220023320223232220022233333223223222222333322322223322232222222222332232323334433333333334545BCCCBCCCBCCBCCBBCCCCBCBBBBBBBBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBABABBABAA9875432220022255555655666667777777787888888888889999998888788875556555355355323344433233235663223333222332232222333333233322223333543333344333333334434432232222202243222023223222022222223323333222223222223220202022222220002222344334433345532222222222222355322200222300332333333220033223433555322223322320220222220330000000220023320223232220022233333223223222222333322322223322232222222222332232323334433333333334545BCCCBCCCBCCBCCBBCCCCBCBBBBBBBBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBABABBABAA98754322200222;
		rom_data[323] <= 3840'h666667777777778888888888999999999888787776566544334333323444443333334552243332323322322223233333333322333333443333333333332335554322222322222233000222343223223233323220222022202222322222022220222202220002223222222233322245202022233344322220222222222322220222233223322332222022332322222232320000200202220024323222232202232222232232222233343333332222323223322222222223332223332334332333333334437BCCBCBCBCBBCBBCCBBBBCBBCBCBCBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBA9886542202222255555556666667777777778888888888999999999888787776566544334333323444443333334552243332323322322223233333333322333333443333333333332335554322222322222233000222343223223233323220222022202222322222022220222202220002223222222233322245202022233344322220222222222322220222233223322332222022332322222232320000200202220024323222232202232222232232222233343333332222323223322222222223332223332334332333333334437BCCBCBCBCBBCBBCCBBBBCBBCBCBCBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBA98865422022222;
		rom_data[324] <= 3840'h666666777777777888888889899999999888788777555543334433333444344433333553253322323322233332323333332232443332444333433333322334575322222322222202202224433020233222332220002222222023553022022222020220222220002022202332222334222202233233022322200233223223322223220220020222222202220222222232222002320220200224223332222223332223232233222233443332332322323222322222022023222232223334333333333333348BCCCCCBCBCCCCCBBCCCCBCBCBBBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBABA987544220222255555555666666777777777888888889899999999888788777555543334433333444344433333553253322323322233332323333332232443332444333433333322334575322222322222202202224433020233222332220002222222023553022022222020220222220002022202332222334222202233233022322200233223223322223220220020222222202220222222232222002320220200224223332222223332223232233222233443332332322323222322222022023222232223334333333333333348BCCCCCBCBCCCCCBBCCCCBCBCBBBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBABA9875442202222;
		rom_data[325] <= 3840'h656667777777778888888888999999998888777777544553324443443324433233245652343323333222233333323345542323542232343333433333323344565222033332200220223322332022220222222202020234220223466430023322222222233232200222222333322222222332222232000202022232322342222233202000233244333220020223232220000202000200222223222222202232332332332222232223322232222322223222223202222222222443333334433333333333348BCCCBCBCCCBBCBBCCBBBCBCBCCCBCBBBBBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA987654322222255555555656667777777778888888888999999998888777777544553324443443324433233245652343323333222233333323345542323542232343333433333323344565222033332200220223322332022220222222202020234220223466430023322222222233232200222222333322222222332222232000202022232322342222233202000233244333220020223232220000202000200222223222222202232332332332222232223322232222322223222223202222222222443333334433333333333348BCCCBCBCCCBBCBBCCBBBCBCBCCCBCBBBBBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA9876543222222;
		rom_data[326] <= 3840'h565667777777777888888889899999999888887776555443336423235533533576355532332432323232343232323334423333444344332323333343543343343232233220220222022222232022222233202200022333220032246530023332022322000232222020222222233222024432000222220020223332223533320223222322332222233322200222220202222320000000232032222232222222222223222202332222322222223322232322223222222322223432333333434333333433349CCBCCCBCBBCCCCBBCBCCBCBCBBCCBBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBABABABAAA98764422222355555555565667777777777888888889899999999888887776555443336423235533533576355532332432323232343232323334423333444344332323333343543343343232233220220222022222232022222233202200022333220032246530023332022322000232222020222222233222024432000222220020223332223533320223222322332222233322200222220202222320000000232032222232222222222223222202332222322222223322232322223222222322223432333333434333333433349CCBCCCBCBBCCCCBBCBCCBCBCBBCCBBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBABABABAAA987644222223;
		rom_data[327] <= 3840'h56666667777777788888888898999999988877777655555433543333853443445435443233244333222232223332322332233232234423223323333334333333223322223202023320223202222022323223332220233322202222222233322022322000022224420202220223322233322020332220020200233233222222333332222222202020020202222332233222342022200002003322222202222232222332220322022232333323322232332222222222223222333332323333433333333335ACCCCCCCCCCCBCBCCBCCBCBCBCBCBBCBBBBCBBCBBBBBBBBBBBBBBBBBBBBBBABBBBBBABAA9876543222225555555556666667777777788888888898999999988877777655555433543333853443445435443233244333222232223332322332233232234423223323333334333333223322223202023320223202222022323223332220233322202222222233322022322000022224420202220223322233322020332220020200233233222222333332222222202020020202222332233222342022200002003322222202222232222332220322022232333323322232332222222222223222333332323333433333333335ACCCCCCCCCCCBCBCCBCCBCBCBCBCBBCBBBBCBBCBBBBBBBBBBBBBBBBBBBBBBABBBBBBABAA987654322222;
		rom_data[328] <= 3840'h55666767777777788888888988999999988887777655556534564233543433333455434325444233322220233322322333232232233332322333332323343333222322233322223222002234302232222002222200233320233222000232222002220000002235422222232222202255300233443023222220022232202222332232222220220000200222333322342202220022200000024422220222223222023322220222220232222223322232323222220222222232223222233233332333333436BCBCBCBCCCCBCBCCBCCBCCCBCBCBCBBBBBBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBABA9987554322225555555555666767777777788888888988999999988887777655556534564233543433333455434325444233322220233322322333232232233332322333332323343333222322233322223222002234302232222002222200233320233222000232222002220000002235422222232222202255300233443023222220022232202222332232222220220000200222333322342202220022200000024422220222223222023322220222220232222223322232323222220222222232223222233233332333333436BCBCBCBCCCCBCBCCBCCBCCCBCBCBCBBBBBBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBABA998755432222;
		rom_data[329] <= 3840'h55656767777777888888888899999999888887777765555534554443434433434434444433343323222322223222223223222343332333323333333223332333322222023320233220222234302232022020220202022202233202002222222222222020202222222023442020222244223223332222222222222222222223222332233223202022222033322222220020000022000000024322223202023222203222222022222222222333222223232322022202222232222322233223332333333447BCCCCCCCBCBCCCBCCBCCBCBCBCBBBBCBCBBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBAAAAAA988754432225555555555656767777777888888888899999999888887777765555534554443434433434434444433343323222322223222223223222343332333323333333223332333322222023320233220222234302232022020220202022202233202002222222222222020202222222023442020222244223223332222222222222222222223222332233223202022222033322222220020000022000000024322223202023222203222222022222222222333222223232322022202222232222322233223332333333447BCCCCCCCBCBCCCBCCBCCBCBCBCBBBBCBCBBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBAAAAAA98875443222;
		rom_data[330] <= 3840'h55666667777777788888888889999999988887777765444433434543433344333343465433332233232222222222322222443355322233332233333323233232332222222222222000233222200022023222022220200000220223200022022222332202320222222233332022022224442202000020022322222224322223222233232222222223222223020200000022200200202002023222222220022222222322223222233222222332222222222222202022222222222222233233433432333347BCCBCCBCCCCBCBCCBCCBCBCBCBCCCBBBBBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA98765432324555555555666667777777788888888889999999988887777765444433434543433344333343465433332233232222222222322222443355322233332233333323233232332222222222222000233222200022023222022220200000220223200022022222332202320222222233332022022224442202000020022322222224322223222233232222222223222223020200000022200200202002023222222220022222222322223222233222222332222222222222202022222222222222233233433432333347BCCBCCBCCCCBCBCCBCCBCBCBCBCCCBBBBBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBA9876543232;
		rom_data[331] <= 3840'h55566667777777888888888889999999988887777765433423433433333344432352357525322222222220222222222223443334323233323333333332323323333223322222200002322202002022223420220222202002300234202022222224554202220243223222220220222235642200000000000022000225322222222233220022233222222202002020202022202002202222022220222220222323223232233222222232222222223222222202222022202223222232333333334432333348BCCCCBCCBCBCCCBCCBCCCCCCBCBBBCCCCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBAA99875433225555555555566667777777888888888889999999988887777765433423433433333344432352357525322222222220222222222223443334323233323333333332323323333223322222200002322202002022223420220222202002300234202022222224554202220243223222220220222235642200000000000022000225322222222233220022233222222202002020202022202002202222022220222220222323223232233222222232222222223222222202222022202223222232333333334432333348BCCCCBCCBCBCCCBCCBCCCCCCBCBBBCCCCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBAA9987543322;
		rom_data[332] <= 3840'h55556667777777778888888888999999988887776765433343433323334454332233245524334222222222222222223223322233433333333333322333233332233323322202202002200000020223233320020222300034430222002022222034444222002022222220222200222234432220002200000223202222022322343334220202223322023200222020222000020002000322022002222022232223233222202223202322222222222222322222222202202322223233333433334332323458CCCBCCCCCCCCBCCCBCBCBBCBCBCCCBBBCBCBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBABBB99875433325455555555556667777777778888888888999999988887776765433343433323334454332233245524334222222222222222223223322233433333333333322333233332233323322202202002200000020223233320020222300034430222002022222034444222002022222220222200222234432220002200000223202222022322343334220202223322023200222020222000020002000322022002222022232223233222202223202322222222222222322222222202202322223233333433334332323458CCCBCCCCCCCCBCCCBCBCBBCBCBCCCBBBCBCBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBABBB9987543332;
		rom_data[333] <= 3840'h5566666777777778888888888989999998887777667545434333443333344433223444442565522222022022222222333222322354343334433333332323323433320222202222222200002200202232020202002222024343220002002220224332220202220020222220200202202222200202222000222322232002202233323433300220222220202332022220000020222020020023222022022232222322222222223222222222222220222233222222222202222222232333343333322323345ACBCBCBCBCBCCCCBCCCCBCCCCBCBBBCCBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABAA987544222545555555566666777777778888888888989999998887777667545434333443333344433223444442565522222022022222222333222322354343334433333332323323433320222202222222200002200202232020202002222024343220002002220224332220202220020222220200202202222200202222000222322232002202233323433300220222220202332022220000020222020020023222022022232222322222222223222222222222220222233222222222202222222232333343333322323345ACBCBCBCBCBCCCCBCCCCBCCCCBCBBBCCBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABAA987544222;
		rom_data[334] <= 3840'h5555666667777778788888888899999998887777667555334333552233543333322344332464320222222222222022333322222354433445433333332332322333330202233322233020022022222020202200002220223222220200002020222220020003322002022022220200200222022320000002002332222202220222022532222222222322020222222220023202020002202222222002022232222222222222222322222222222020220232222202220222322222223333233333323233345ACCCCCCCCCCBCBCBCBCBCCBCBCCCCCBBBBCBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBABBBBABBBA9887553322455555555555666667777778788888888899999998887777667555334333552233543333322344332464320222222222222022333322222354433445433333332332322333330202233322233020022022222020202200002220223222220200002020222220020003322002022022220200200222022320000002002332222202220222022532222222222322020222222220023202020002202222222002022232222222222222222322222222222020220232222202220222322222223333233333323233345ACCCCCCCCCCBCBCBCBCBCCBCBCCCCCBBBBCBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBABBBBABBBA9887553322;
		rom_data[335] <= 3840'h5556666677777777888888888889999988887776677654334323443323543542322433432343222220222220222222333322222334444444433232323433223333233222033432232220220002222203202220022220222220222000222022320202000022220020020024320200222002020200000020020332200223200222203332033220222222322002220002332000220002022223322200222222222233322220222222222002222022222222222223532222223322333333333333223233347BCCBCCCCBCBCCCCCCCCBCBCCCBCBCBCBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBAA9987543222454555555556666677777777888888888889999988887776677654334323443323543542322433432343222220222220222222333322222334444444433232323433223333233222033432232220220002222203202220022220222220222000222022320202000022220020020024320200222002020200000020020332200223200222203332033220222222322002220002332000220002022223322200222222222233322220222222222002222022222222222223532222223322333333333333223233347BCCBCCCCBCBCCCCCCCCBCBCCCBCBCBCBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBAA9987543222;
		rom_data[336] <= 3840'h5555666667777777788888888898999998887766567644453333343323433432233332245444222222022022222222332222234434344443443333333322222232323323222322233220202020222202220222223220222020202222222202220020033202002200000222200023320200000000000020022022220220022352222222222202233302202023222002320002220022220223220220002222222333222222222322222222203223222222202025622222222222233332333323222333348BCBCBCBCCCCCCCCBCBCCBCBCBCBCCCCBBBBCBCBCBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBAA8886543222454555555555666667777777788888888898999998887766567644453333343323433432233332245444222222022022222222332222234434344443443333333322222232323323222322233220202020222202220222223220222020202222222202220020033202002200000222200023320200000000000020022022220220022352222222222202233302202023222002320002220022220223220220002222222333222222222322222222203223222222202025622222222222233332333323222333348BCBCBCBCCCCCCCCBCBCCBCBCBCBCCCCBBBBCBCBCBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBAA8886543222;
		rom_data[337] <= 3840'h5555666677777777878888888889999998887765557644563433333343323332343332258543222222322202220222344323334433444554444333223232222323333332322222022202202220022002330022220202222200202222200202022222222020000202232202022233322022220002200020000023223222202233222222200003332222022220222022200022200222022222202200222232023333222222223223222220202222322220200224220222222222233333333332223323349CCCCBCCCCCCCBCCCCCCBCBCBCCCBCBCCCCCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBABBBBBA98876543202445455555555666677777777878888888889999998887765557644563433333343323332343332258543222222322202220222344323334433444554444333223232222323333332322222022202202220022002330022220202222200202222200202022222222020000202232202022233322022220002200020000023223222202233222222200003332222022220222022200022200222022222202200222232023333222222223223222220202222322220200224220222222222233333333332223323349CCCCBCCCCCCCBCCCCCCBCBCBCCCBCBCCCCCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBABBBBBA98876543202;
		rom_data[338] <= 3840'h555555666777777778888888888989999888775555774454343443334333333334223235543302222222222022220223433232332334444434553323233222323333343232200222020200002200022222220200002222022222222200002022422223300202002234322022322222222220000022002000202222222220000222220000002343222222222202222222000200002002022222222202022222453322222220222322222222202232222202022220222222223322233333333223232335BCCBCCCBCBCCCCBCBCBCCCCCCCBBCBCBBCBCBCBCBCBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBAA9887553222044455555555555666777777778888888888989999888775555774454343443334333333334223235543302222222222022220223433232332334444434553323233222323333343232200222020200002200022222220200002222022222222200002022422223300202002234322022322222222220000022002000202222222220000222220000002343222222222202222222000200002002022222222202022222453322222220222322222222202232222202022220222222223322233333333223232335BCCBCCCBCBCCCCBCBCBCCCCCCCBBCBCBBCBCBCBCBCBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBAA98875532220;
		rom_data[339] <= 3840'h555556667777777778888888889899988887665555775333333433543444323554223333443322222220220220202223332222232344434335553233232222223332333453202202020020020002022200222022232322222202220002000222220023223420002223202022320022222200232222020000022202000022220000200020222233323322222222220020000000020202022202022000000222552222222222222222222222222222222220202202032222223323333233332232322335BCCCCBCCCCCBCCBCCCCCBBCBBCCCBBCBCCCBCBCBCBBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBAA99876543200044545555555556667777777778888888889899988887665555775333333433543444323554223333443322222220220220202223332222232344434335553233232222223332333453202202020020020002022200222022232322222202220002000222220023223420002223202022320022222200232222020000022202000022220000200020222233323322222222220020000000020202022202022000000222552222222222222222222222222222222220202202032222223323333233332232322335BCCCCBCCCCCBCCBCCCCCBBCBBCCCBBCBCCCBCBCBCBBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBAA998765432000;
		rom_data[340] <= 3840'h555565666677777777888888889899898877655554575433343334553445434553223333554344222220222222022233222222023334433434544233232223322333333453232220200220200022022002322222223222222200002022020020000000225520000202002322022000222002332202002000022222300002222202020022020223222322222202220200020002000020000202222220220203332222022222322222222222022222222222020220223202223322332333332233222337BCCBCCCCCBCCCBCBCBCBCCBCCCBBCCBCBCBCBCBCBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBA98875442222044445555555565666677777777888888889899898877655554575433343334553445434553223333554344222220222222022233222222023334433434544233232223322333333453232220200220200022022002322222223222222200002022020020000000225520000202002322022000222002332202002000022222300002222202020022020223222322222202220200020002000020000202222220220203332222022222322222222222022222222222020220223202223322332333332233222337BCCBCCCCCBCCCBCBCBCBCCBCCCBBCCBCBCBCBCBCBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBA988754422220;
		rom_data[341] <= 3840'h555556666777777787888888888998888877655544555444343345533335323443223334675334322220220220200222222202232024433444333222332234223223332333333422002232200222000220222020220003320200020222220202000000024420002200023320202020200020222000020222222323200200020202200222202232222222222220000002022022020220022020202022222202322222222202220222322220222023222222020200222222233223322333333222233349CCCCCBCBCCCBCCBCCCCCBCCBCBCCBBCBCCCBCBCBCBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBAA88765432200044455455555556666777777787888888888998888877655544555444343345533335323443223334675334322220220220200222222202232024433444333222332234223223332333333422002232200222000220222020220003320200020222220202000000024420002200023320202020200020222000020222222323200200020202200222202232222222222220000002022022020220022020202022222202322222222202220222322220222023222222020200222222233223322333333222233349CCCCCBCBCCCBCCBCCCCCBCCBCBCCBBCBCCCBCBCBCBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBAA887654322000;
		rom_data[342] <= 3840'h55555566667777777778888888898988887755555445444433354332333333333223323456432222222222222022022223232232222243344433322334332333223333322222220202222000022022023232002302000220200222022033222000000000220000002233200022020202200000000020200222222222200202022220232002222320220202020020202000000220000002200020222202222222022022220222022224222022222322220202222222222233322223223333222322345BCCCCCCCCCBCCCCCCCCCCCBCCBCCBCCBCBCBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBA98775543220004444455555555566667777777778888888898988887755555445444433354332333333333223323456432222222222222022022223232232222243344433322334332333223333322222220202222000022022023232002302000220200222022033222000000000220000002233200022020202200000000020200222222222200202022220232002222320220202020020202000000220000002200020222202222222022022220222022224222022222322220202222222222233322223223333222322345BCCCCCCCCCBCCCCCCCCCCCBCCBCCBCCBCBCBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBA9877554322000;
		rom_data[343] <= 3840'h55555566666777777788888888898988877655544345533333244332343323433233223333332222022020202202022233222322222333333333333334422223323332200002200002000000200023232320222022023222200222202222202220000222000002222233202222332222320000002000000000022322020022222222202223222200222320200022000200000000222222000220002020222222022222220222220234322202223332322022020222222332222222233333223222347CCCCCCBCBCCCBCBCCBCBCCCCCCBCBCBCBCCCBCBCBCBCBBCBBBCBBBBBBBBBBBBBBBBBBBBBAA98765432200204445455555555566666777777788888888898988877655544345533333244332343323433233223333332222022020202202022233222322222333333333333334422223323332200002200002000000200023232320222022023222200222202222202220000222000002222233202222332222320000002000000000022322020022222222202223222200222320200022000200000000222222000220002020222222022222220222220234322202223332322022020222222332222222233333223222347CCCCCCBCBCCCBCBCCBCBCCCCCCBCBCBCBCCCBCBCBCBCBBCBBBCBBBBBBBBBBBBBBBBBBBBBAA9876543220020;
		rom_data[344] <= 3840'h55555556666777777778888888898888777655444445533333244433333333333243322233322022222222022222222233223322233443333332432334332222222222222220000200222000002223202202222202232220202022220202202022002332000222220000000233442222220000202000200000023320020000220233222222020222022202202222000002000202202020200022202220222220022222222222222234320220223442202222222222222222222022233333222222349CCCCCCCCCCBCCCCBCCCCBCCBCBCBCBBCBCBCBCBCBCBCCCBBCBBBBBBBBBBBBBBBBBBBBBBBB988755432020004444454555555556666777777778888888898888777655444445533333244433333333333243322233322022222222022222222233223322233443333332432334332222222222222220000200222000002223202202222202232220202022220202202022002332000222220000000233442222220000202000200000023320020000220233222222020222022202202222000002000202202020200022202220222220022222222222222234320220223442202222222222222222222022233333222222349CCCCCCCCCCBCCCCBCCCCBCCBCBCBCBBCBCBCBCBCBCBCCCBBCBBBBBBBBBBBBBBBBBBBBBBBB98875543202000;
		rom_data[345] <= 3840'h5555556666677777788888888888888777655444343554333323443433333443333222234233322222222222222055323223233333334433333232223432232222222222220202222222000022232222022222222232222200222222222022220220222000222002202200222332222200000000002202200202202022200220222202020020222202022002220002202000022000002220020202222232222022232222222220223322220222333220223203222222222222022233333422222235ACCCCCCCCCCCCBCCCCBCCCCBCCCCCBCBCBCBCBCBCBCBCBBBCBBCBCBBBBBBBBBBBBBBBBBAAA98775533220000444454555555556666677777788888888888888777655444343554333323443433333443333222234233322222222222222055323223233333334433333232223432232222222222220202222222000022232222022222222232222200222222222022220220222000222002202200222332222200000000002202200202202022200220222202020020222202022002220002202000022000002220020202222232222022232222222220223322220222333220223203222222222222022233333422222235ACCCCCCCCCCCCBCCCCBCCCCBCCCCCBCBCBCBCBCBCBCBCBBBCBBCBCBBBBBBBBBBBBBBBBBAAA98775533220000;
		rom_data[346] <= 3840'h5555555666677777777888888888887776555443433455333323333442244433222232345223322222202222002255320223322332333333333222222322222222202020220002222222000222220202022222202223220020222222222200000022000002020022222200022220002000202000000000222220200022020202000022022200022200202022202022020000202220000220000202330220222222254202220202222222222222232222222222222222222022222233234422232236CCCCCCBCBCBCCCBCBCCBCBCCCCBCBCBCBCBCBCBCBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBAA998765432202000444454455555555666677777777888888888887776555443433455333323333442244433222232345223322222202222002255320223322332333333333222222322222222202020220002222222000222220202022222202223220020222222222200000022000002020022222200022220002000202000000000222220200022020202000022022200022200202022202022020000202220000220000202330220222222254202220202222222222222232222222222222222222022222233234422232236CCCCCCBCBCBCCCBCBCCBCBCCCCBCBCBCBCBCBCBCBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBAA998765432202000;
		rom_data[347] <= 3840'h5555555666777777778888888888887775554434333455543333333442244323223322333233222220222020020224322022332223333333432222223332222222222222000200020222000202202222202220022022200022222220220002000202000220200022222002002022002022022200000000020220202222200202200202022202002000220220020022200002220200022200202222220002202220253220020202222202020222222222202222222222222222233233334322222348CCCCCCCCCCCCCBCCCCCCCCCBCBCBCBCBCBCBCBCBCBCBCBCBBCBCBBCBBBBBBBBBBBBBBBAA9987755332220000344444545555555666777777778888888888887775554434333455543333333442244323223322333233222220222020020224322022332223333333432222223332222222222222000200020222000202202222202220022022200022222220220002000202000220200022222002002022002022022200000000020220202222200202200202022202002000220220020022200002220200022200202222220002202220253220020202222202020222222222202222222222222222233233334322222348CCCCCCCCCCCCCBCCCCCCCCCBCBCBCBCBCBCBCBCBCBCBCBCBBCBCBBCBBBBBBBBBBBBBBBAA9987755332220000;
		rom_data[348] <= 3840'h555555556667777778788888888887766555443434334555433323443233333232332233233332222202222220200323222222332233433343222322335423222224554220220200022022020200232220022002222202200200202202200000220002022000020022220020000220200020220020000000222222023220022222200202002200000222222222200000000232220002222220022222202222222222202022202022222202202022202020200222022222222223223233320222225ACCCCCCCBCCCCCCCCCCBCCBCCCCCCCCBCBCBCBCBCBCBCBCBCCBBBCBBBBBBBBBBBBBBBBBA9988765432220020044444445555555556667777778788888888887766555443434334555433323443233333232332233233332222202222220200323222222332233433343222322335423222224554220220200022022020200232220022002222202200200202202200000220002022000020022220020000220200020220020000000222222023220022222200202002200000222222222200000000232220002222220022222202222222222202022202022222202202022202020200222022222222223223233320222225ACCCCCCCBCCCCCCCCCCBCCBCCCCCCCCBCBCBCBCBCBCBCBCBCCBBBCBBBBBBBBBBBBBBBBBA99887654322200200;
		rom_data[349] <= 3840'h555555566666777777788888888877765554443433334554343223332234322222222353223322232222202222222223320222232233334433222232234532322024653322202022220233322002202202020023320002000002222020022020220222020000322222000020002222000002220000002020222020023220022222002022000022022222220222020220000233220022322020222322020022202222202220020220222022022222202200202202222222220223223332222222235BCCCCCCCCCCCCCBCBCBCCCCCBCCBBCBCBCBCBCBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBAAA9887654432200200043444454555555566666777777788888888877765554443433334554343223332234322222222353223322232222202222222223320222232233334433222232234532322024653322202022220233322002202202020023320002000002222020022020220222020000322222000020002222000002220000002020222020023220022222002022000022022222220222020220000233220022322020222322020022202222202220020220222022022222202200202202222222220223223332222222235BCCCCCCCCCCCCCBCBCBCCCCCBCCBBCBCBCBCBCBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBAAA98876544322002000;
		rom_data[350] <= 3840'h555555555666677777878888888777755554443334344554333323232343322332222443233222232222222220220222222223222333333332222322222322222222223220000022220233220022000002222002220022020022200200230000020000022000344302200020002002220002000000000000020202202200002000222220222002022022220222202000200222200002220002023322200222202222022022202222222200202220220202020202223222222222322323202222237CCCCCBCBCCCCBCCCCCCCBCBCCCCCBCBCBCBCBCBCBCBCBCBCCBCBBBBCBBBBBBBBBBBBAAA99876554322020000034444444555555555666677777878888888777755554443334344554333323232343322332222443233222232222222220220222222223222333333332222322222322222222223220000022220233220022000002222002220022020022200200230000020000022000344302200020002002220002000000000000020202202200002000222220222002022022220222202000200222200002220002023322200222202222022022202222222200202220220202020202223222222222322323202222237CCCCCBCBCCCCBCCCCCCCBCBCCCCCBCBCBCBCBCBCBCBCBCBCCBCBBBBCBBBBBBBBBBBBAAA998765543220200000;
		rom_data[351] <= 3840'h455555556566777777788888888776655554434443445544444322333322322332223322243323432222002222002220202332223332442332322232222222223220022322022222022000000022000222220020202202222022000022200000222000000020020002000220000020222200000000000002200220022000020222034202022000000023322222202000002022000002220000035322002222022220220222222024420022020222202202002202222222220232323232222202259CCCBCCCCCCCCCCBCCBCCCCCCBCBCCBCBCBBCBBCBCBCBCBCBBCBBCBCBBBBBBBBBBBBAAA988776543322000000034344445455555556566777777788888888776655554434443445544444322333322322332223322243323432222002222002220202332223332442332322232222222223220022322022222022000000022000222220020202202222022000022200000222000000020020002000220000020222200000000000002200220022000020222034202022000000023322222202000002022000002220000035322002222022220220222222024420022020222202202002202222222220232323232222202259CCCBCCCCCCCCCCBCCBCCCCCCBCBCCBCBCBBCBBCBCBCBCBCBBCBBCBCBBBBBBBBBBBBAAA9887765433220000000;
		rom_data[352] <= 3840'h45555555666677777777888888877655555444444445554344333223232233223233322223322332222220202222022222223332233332333323222222222203532020222202200020000200000000002200220200020023322020220000002202000002000000000000022000000002020000000000020220222022200000222222200202022002023430243200020002000020000232200023443222223222020202222222023442020022202020020002020022222222332322332220222225ACCCCBCCCCCCCBCCBCCCBCCBCCCCCBCCBCCBBBBCBCBCBCBCCBCBBBBBBBBBBBBBBBBAA9998876544322202000004344444545555555666677777777888888877655555444444445554344333223232233223233322223322332222220202222022222223332233332333323222222222203532020222202200020000200000000002200220200020023322020220000002202000002000000000000022000000002020000000000020220222022200000222222200202022002023430243200020002000020000232200023443222223222020202222222023442020022202020020002020022222222332322332220222225ACCCCBCCCCCCCBCCBCCCBCCBCCCCCBCCBCCBBBBCBCBCBCBCCBCBBBBBBBBBBBBBBBBAA999887654432220200000;
		rom_data[353] <= 3840'h45555555566667777778888887776655555554545555555334432332333233322332322322232332022222020222222222223332233323332332222220222222342222202222000000020000200020202020220022020202320002200000000200220220220000000000200000002220202200000000000002000022202023322200002000000220202222232202000220020020202232000222332222343222222202222020022220220222220202020220202222222222222223323222222237BCCBCCCBCCCCCCCCCCBCCCCCCBCBCCBCBCBCCBBCBCBCBCBBBCBBCBCBBCBBBBBBABAA99987765443222200000003443444545555555566667777778888887776655555554545555555334432332333233322332322322232332022222020222222222223332233323332332222220222222342222202222000000020000200020202020220022020202320002200000000200220220220000000000200000002220202200000000000002000022202023322200002000000220202222232202000220020020202232000222332222343222222202222020022220220222220202020220202222222222222223323222222237BCCBCCCBCCCCCCCCCCBCCCCCCBCBCCBCBCBCCBBCBCBCBCBBBCBBCBCBBCBBBBBBABAA9998776544322220000000;
		rom_data[354] <= 3840'h45555555566667777787888877776665555555555555675333323223332233322223223322243322222202222222023222222323323222232323322022222202222222023220200202202220020002220202202202220002020000222000000200000220020000000000000000002022000020000000000002002020200022333200000200000200000020020200000002020002002322200222222222332222222222222022002220002222202202002020202222222222222222333202222349CCCCCBCCBCCCCBCCBCCCCBCBCCBBCBCBCBCBCBCBCBCBCBCBBBCBBBBBBBBBAAABAAA999887654433222020000004344444545555555566667777787888877776665555555555555675333323223332233322223223322243322222202222222023222222323323222232323322022222202222222023220200202202220020002220202202202220002020000222000000200000220020000000000000000002022000020000000000002002020200022333200000200000200000020020200000002020002002322200222222222332222222222222022002220002222202202002020202222222222222222333202222349CCCCCBCCBCCCCBCCBCCCCBCBCCBBCBCBCBCBCBCBCBCBCBCBBBCBBBBBBBBBAAABAAA99988765443322202000000;
		rom_data[355] <= 3840'h5555555566666777777788877777665655555555566777633333232322223332233322333223222223432202202222222222332332322223323323222220202202222002220020020202220002020000200002022022002222020002000000020200000020000000000000200222203200002000000000022000202002222223322220002002220002022022020000002002020002232202222202202222222222322222222202222020222022202202202022222222222222222232322202226BCCCBCCCBCCCCCCCCCCBCCCCCCBCBCBCCBCBBCBBCBCBCBCBBCBBBBBBBBABAAAAAA9998887655433220200000000343444445555555566666777777788877777665655555555566777633333232322223332233322333223222223432202202222222222332332322223323323222220202202222002220020020202220002020000200002022022002222020002000000020200000020000000000000200222203200002000000000022000202002222223322220002002220002022022020000002002020002232202222202202222222222322222222202222020222022202202202022222222222222222232322202226BCCCBCCCBCCCCCCCCCCBCCCCCCBCBCBCCBCBBCBBCBCBCBCBBCBBBBBBBBABAAAAAA9998887655433220200000000;
		rom_data[356] <= 3840'h4455555655667777777788787777766666565556677778743232332232222322343332222344222322532220220020222222222222322244233323202022222302332002222222023322222022200000022002202000000220202200000000222002000000000000002000000343224430000000000000022202002222202222222020020200202220020022020020200200220002322202222020200022202222332322202202020222000220220200220202222220222222232232220222328CCBCCCBCCCCCCCBCBCCCCCCCBCCCBCCCBCBCBCBBBCBCBCBCBBCBBBBBBBAAA9AA999988876554332220020000000334344444455555655667777777788787777766666565556677778743232332232222322343332222344222322532220220020222222222222322244233323202022222302332002222222023322222022200000022002202000000220202200000000222002000000000000002000000343224430000000000000022202002222202222222020020200202220020022020020200200220002322202222020200022202222332322202202020222000220220200220202222220222222232232220222328CCBCCCBCCCCCCCBCBCCCCCCCBCCCBCCCBCBCBCBBBCBCBCBCBBCBBBBBBBAAA9AA999988876554332220020000000;
		rom_data[357] <= 3840'h4555555556667777777788877777666666666667777788853232323332322432233322332345322322323202202220244222222002222463232233222222223322230222002320223320220222000002220020222000000020222200022000022220000000000000022000020232224430200000000222000020002332202020202000000022200320000220200000002000020002222022222220200220222222443220220022020000020222202002020222222222202222332332202202339CCCCCBCCCCCCCCCBCCCBCBCCCBCBCBBBCCBCBCBCCBCBCBCBBBBBBBABAAAAA999988887765543322200200000000434444444555555556667777777788877777666666666667777788853232323332322432233322332345322322323202202220244222222002222463232233222222223322230222002320223320220222000002220020222000000020222200022000022220000000000000022000020232224430200000000222000020002332202020202000000022200320000220200000002000020002222022222220200220222222443220220022020000020222202002020222222222202222332332202202339CCCCCBCCCCCCCCCBCCCBCBCCCBCBCBBBCCBCBCBCCBCBCBCBBBBBBBABAAAAA999988887765543322200200000000;
		rom_data[358] <= 3840'h445555555666677777787888777777776777777777888887432333233332245222333323222432232222220202200223432200222002334333323222222220222022202022222220200232200020020000000000220002022202000002200000002202200002220000000220202002232232000020000002200020333200022022220020020200000002020000000000202000002233020202020202020202223343202020222200200200000200220202022232222222332232223202222226BCCCCCCCCCCCCCCBCCCCCBCCBCCBCCCCBCBBCBCBBCBCBCBCBCBBBBBAAAAA9998888877765543322202000000000033434444445555555666677777787888777777776777777777888887432333233332245222333323222432232222220202200223432200222002334333323222222220222022202022222220200232200020020000000000220002022202000002200000002202200002220000000220202002232232000020000002200020333200022022220020020200000002020000000000202000002233020202020202020202223343202020222200200200000200220202022232222222332232223202222226BCCCCCCCCCCCCCCBCCCCCBCCBCCBCCCCBCBBCBCBBCBCBCBCBCBBBBBAAAAA99988888777655433222020000000000;
		rom_data[359] <= 3840'h555555555666777777778887777777777777777888888998532332333322244222323323233322233222222022022022332222222022223322223232222222022000222222000220000232002222000020000000000000200200020000000000020020000022200000000200000002220220000020000000002020222020022200020002200002000200002020002000222200002242202222222000020202222332220202202022000000200200002020202222222223322222243220022339CCCBCCBCCCCBCBCCBCCCBCCCCCBCCBBCBCCBBCBBBCBCBCBCBBBBBAAA99998888887777655433322020000000000043434444555555555666777777778887777777777777777888888998532332333322244222323323233322233222222022022022332222222022223322223232222222022000222222000220000232002222000020000000000000200200020000000000020020000022200000000200000002220220000020000000002020222020022200020002200002000200002020002000222200002242202222222000020202222332220202202022000000200200002020202222222223322222243220022339CCCBCCBCCCCBCBCCBCCCBCCCCCBCCBBCBCCBBCBBBCBCBCBCBBBBBAAA999988888877776554333220200000000000;
		rom_data[360] <= 3840'h44555555556667777777787888777777777878888889999853233323333223322222232223222233220202020200022022002222202232232222232322222320222022022222002000022220200000002022200020000000200000220000000000220222330000002022002022200002000000000000222020200002022200002000002222000023200020202000000022220000023202002020202020202222222222200202220202000000002000020222222220222332222233220202235ACCCCCCCBCCCCCCBCCCCCCCCBCCCCBCCBCBCBCBCBCBCBBCCBBBBAAA999988888887776655443222020000000000003434444444555555556667777777787888777777777878888889999853233323333223322222232223222233220202020200022022002222202232232222232322222320222022022222002000022220200000002022200020000000200000220000000000220222330000002022002022200002000000000000222020200002022200002000002222000023200020202000000022220000023202002020202020202222222222200202220202000000002000020222222220222332222233220202235ACCCCCCCBCCCCCCBCCCCCCCCBCCCCBCCBCBCBCBCBCBCBBCCBBBBAAA99998888888777665544322202000000000000;
		rom_data[361] <= 3840'h5555555556667777777788888887778788888888899999A973233222332233322233232222222332222220200002220200202422222222222222222222222222220220002202000222202020002000200022000020232000200002200020000020020223432000000220222200000020000002000000000020200000202000020002222200220202020222000002000020202020223202000202022200222223323222200002022220000000020020200002222332223222222233220222338CCCCCBCCCCBCCBCCCBCBCCBCCCBCBCBCBCBCBCBCBCBBBCBCBBBAA9999888887777765555443222200000000000000343444445555555556667777777788888887778788888888899999A973233222332233322233232222222332222220200002220200202422222222222222222222222222220220002202000222202020002000200022000020232000200002200020000020020223432000000220222200000020000002000000000020200000202000020002222200220202020222000002000020202020223202000202022200222223323222200002022220000000020020200002222332223222222233220222338CCCCCBCCCCBCCBCCCBCBCCBCCCBCBCBCBCBCBCBCBCBBBCBCBBBAA9999888887777765555443222200000000000000;
		rom_data[362] <= 3840'h45555555556667777777888787888888888888888999999A84333322333233233332222022222322202020202020020222022320222222222222202020222220220000020002200202000002000002020000200000220000000000002202000222000002432000000000022200000222000000000000000020000000220200002000220222023300002002000000000000202200222000002202000222222222222222220220223302020202000020332220222220232222222232020202349CCCBCCBCBCCBCCCBCCCCBCCCBCCBCCBCBCBCBCBCBCBBBCBBBABA998888877777765555443332202000000000000003343444445555555556667777777888787888888888888888999999A84333322333233233332222022222322202020202020020222022320222222222222202020222220220000020002200202000002000002020000200000220000000000002202000222000002432000000000022200000222000000000000000020000000220200002000220222023300002002000000000000202200222000002202000222222222222222220220223302020202000020332220222220232222222232020202349CCCBCCBCBCCBCCCBCCCCBCCCBCCBCCBCBCBCBCBCBCBBBCBBBABA99888887777776555544333220200000000000000;
		rom_data[363] <= 3840'h55555555566677777777888888888888888888999999AAAA9533332333233222233322222222222222202020000020202222222220022222222222220223320202000020002020200000000200000020000000002200000200000000020222220002000232200000002002002020002020020200000000020000000022200202200000222002330222002020000000002000200022202022022002202222200222222200222222322020200200000222202202202022223222232220202236BCCCCCCCCCCCCCBCCCBCCCCBCCCCCBBCCBCBCBCBCBCBCBBCBBAA9988877776665555554433322200000000000000003434444455555555566677777777888888888888888888999999AAAA9533332333233222233322222222222222202020000020202222222220022222222222220223320202000020002020200000000200000020000000002200000200000000020222220002000232200000002002002020002020020200000000020000000022200202200000222002330222002020000000002000200022202022022002202222200222222200222222322020200200000222202202202022223222232220202236BCCCCCCCCCCCCCBCCCBCCCCBCCCCCBBCCBCBCBCBCBCBCBBCBBAA998887777666555555443332220000000000000000;
		rom_data[364] <= 3840'h455555555667677777877888888888888888999999A9AAAAA743333333243222322322222222222222200202202002222022202022022222220220222023320200000222000220202022002220002000000000202220000002220000020020202002000020000200002000020002000002200000000002002000200002022000020000022002220002002020200200202000000222220020200020202222222022222222020222222000002022020220220020220202242223232222022348CCCCCCBCCCBCBCCCBCCCCBCCCCBCBCCBCBCBCBCBCBCBBBBBBAA998877765555555554443322220200000000000000043444444455555555667677777877888888888888888999999A9AAAAA743333333243222322322222222222222200202202002222022202022022222220220222023320200000222000220202022002220002000000000202220000002220000020020202002000020000200002000020002000002200000000002002000200002022000020000022002220002002020200200202000000222220020200020202222222022222222020222222000002022020220220020220202242223232222022348CCCCCCBCCCBCBCCCBCCCCBCCCCBCBCCBCBCBCBCBCBCBBBBBBAA9988777655555555544433222202000000000000000;
		rom_data[365] <= 3840'h455555556666777777788888888888888899999AAAAAAAAAB84323232233332232232233232222222020202000020222222202222002222220222222022222222000000200220022200222020000000002000020232000000020200202020002202000000000000000000020020202022000000000000000000220002022000020222022000220022002020000000000000000202220020200202202202022220220202020020222020202002020200200222022220233222222320022235BCCCCBCCCBCCCCCBCBCBCCCCBCCCCCBBCCCCCBCBBCBCBCBBBAA9888766555555444443333232200000000000000000034344445455555556666777777788888888888888899999AAAAAAAAAB84323232233332232232233232222222020202000020222222202222002222220222222022222222000000200220022200222020000000002000020232000000020200202020002202000000000000000000020020202022000000000000000000220002022000020222022000220022002020000000000000000202220020200202202202022220220202020020222020202002020200200222022220233222222320022235BCCCCBCCCBCCCCCBCBCBCCCCBCCCCCBBCCCCCBCBBCBCBCBBBAA98887665555554444433332322000000000000000000;
		rom_data[366] <= 3840'h555555555666777777788888888888899999A9A9AAAAAAAAA95322323223323232222223232222222222202022002002322200220222222222222222202000233200200200002002020223202000000020000002222222020000022222220200020000000000000000020220220020222022000000000000000000020002202200020022002222020000020220000020000020002220200002020000222022002020200220000002020200200220020020202020222233202222200022238CCCCCCCBCCCCCBCCCCCCBCBCCCCCCBCCBCBBCBCBBCBCBBBAA998887655544444444333232222020000000000000000034344444555555555666777777788888888888899999A9A9AAAAAAAAA95322323223323232222223232222222222202022002002322200220222222222222222202000233200200200002002020223202000000020000002222222020000022222220200020000000000000000020220220020222022000000000000000000020002202200020022002222020000020220000020000020002220200002020000222022002020200220000002020200200220020020202020222233202222200022238CCCCCCCBCCCCCBCCCCCCBCBCCCCCCBCCBCBBCBCBBCBCBBBAA9988876555444444443332322220200000000000000000;
		rom_data[367] <= 3840'h5555555566676777788788888888898999999A9AAAAAAAAAAB733323323233222223322222322223322002202020022222022202002222234222200202022022202200000022002002223320002000000200000022222000202000022020220020020000000000020002020200002020222000000000020000200200022000002020000000002000000000202000000020000000222200220222022020020020200220220202202002202000000000202220220220223222222220222225ACCBCBCCCCBCBCCCBBCBCCCCCBCBCBCBCCCCCBCBBCCBCBABA99887765444343333333322222202000000000000000000343444455555555566676777788788888888898999999A9AAAAAAAAAAB733323323233222223322222322223322002202020022222022202002222234222200202022022202200000022002002223320002000000200000022222000202000022020220020020000000000020002020200002020222000000000020000200200022000002020000000002000000000202000000020000000222200220222022020020020200220220202202002202000000000202220220220223222222220222225ACCBCBCCCCBCBCCCBBCBCCCCCBCBCBCBCCCCCBCBBCCBCBABA99887765444343333333322222202000000000000000000;
		rom_data[368] <= 3840'h455555556666777777788888888898999999A9A9AAAAAAAAAB842333323233322223222232222222220202220200202222200000200222222322220220200200020000000202202002222200000000200002000022202002220000000202202022000000000000002202200002200000200000000000020000000200002000002000222000000000000000220000000020020002222020020202020200202020222220222020202002200200020200202202022022222222222220022237CCCBCCBCCCCCCCCBCCCCCCCBCCCCBCCCBCBBBCBCCBBBBAAAA9887755444333332332222222020020000000000000000043444454455555556666777777788888888898999999A9A9AAAAAAAAAB842333323233322223222232222222220202220200202222200000200222222322220220200200020000000202202002222200000000200002000022202002220000000202202022000000000000002202200002200000200000000000020000000200002000002000222000000000000000220000000020020002222020020202020200202020222220222020202002200200020200202202022022222222222220022237CCCBCCBCCCCCCCCBCCCCCCCBCCCCBCCCBCBBBCBCCBBBBAAAA98877554443333323322222220200200000000000000000;
		rom_data[369] <= 3840'h55555556666677777788888888888999999A9A9AAAAAAAAAAB95333332333332222222222222220222220232002020220222002222000202332002020200000202020202022200000002002200000000020000000002200020000000002020222220000000000000000200022200002000000000000000000000000000000000020000000000200200000200002000000000002230000220000202000220002222020200220222022020000000000002002202022220222222220222324ACCCCCCCCCBCBCCBCCCCCBCCCCBCBCBCBCBCCBBBBBBBBAAA99887755543322222222222220202000000000000000000003444444555555556666677777788888888888999999A9A9AAAAAAAAAAB95333332333332222222222222220222220232002020220222002222000202332002020200000202020202022200000002002200000000020000000002200020000000002020222220000000000000000200022200002000000000000000000000000000000000020000000000200200000200002000000000002230000220000202000220002222020200220222022020000000000002002202022220222222220222324ACCCCCCCCCBCBCCBCCCCCBCCCCBCBCBCBCBCCBBBBBBBBAAA9988775554332222222222222020200000000000000000000;
		rom_data[370] <= 3840'h555555566666777777888888888888899999A9A9AAAAAAAAABA6423333232232222222222222222202202232020022022022220020200022222200002020000000022202202022020000000000220000000000020200000232000000000220002200000000002200020020202220200000000000000000202000000000000200002200000000000000000200002000000000000322000020022202200000220222022220002022022220000020000202000222022222202223222232227CCCBBCBCCCCCCBCCCBCBCCBCBCCCCCCBCCCCBBCBCBCBAA99987766544322222222022020002002000000000000000000034344444555555566666777777888888888888899999A9A9AAAAAAAAABA6423333232232222222222222222202202232020022022022220020200022222200002020000000022202202022020000000000220000000000020200000232000000000220002200000000002200020020202220200000000000000000202000000000000200002200000000000000000200002000000000000322000020022202200000220222022220002022022220000020000202000222022222202223222232227CCCBBCBCCCCCCBCCCBCBCCBCBCCCCCCBCCCCBBCBCBCBAA999877665443222222220220200020020000000000000000000;
		rom_data[371] <= 3840'h55555556666777777788888888888999999A9A9AAAAAAAAAAAB953334222222222222220222222222220222200020222222220022002002020020000020000002000000020220002000020000002000002200000000002222000000022020022200000000000000000220002220022000000000000000000000000000000000200020200000000000000020000000000000000222000000022322200002202220222020020222022220000000002000202020022222022222222223224ACCCCCCCCBCCBCCBCBCCCCCCCCBCBBCBCBBBCBCBBBBBAA99887765543322220202020000000002000000000000000000004444445555555556666777777788888888888999999A9A9AAAAAAAAAAAB953334222222222222220222222222220222200020222222220022002002020020000020000002000000020220002000020000002000002200000000002222000000022020022200000000000000000220002220022000000000000000000000000000000000200020200000000000000020000000000000000222000000022322200002202220222020020222022220000000002000202020022222022222222223224ACCCCCCCCBCCBCCBCBCCCCCCCCBCBBCBCBBBCBCBBBBBAA9988776554332222020202000000000200000000000000000000;
		rom_data[372] <= 3840'h55555565666777777777888888889899999999A9AAAAAAAAAABB73234323232222222222222222222222002220200022222202002000202222202000000000000200000022220200000000000000000000202002020002200000000222200020200002000000000000000200220022000000000000002000000200000020002002000020000000000000202000000200000000222202020023320000022022222002000020022020222000000000000202020222222202222222223237CCCCCCCBCCBCCCBCCCCCBCBCCCCCCBCCBCCBCCBBBBBAA998877555433220200000000000000000000000000000000000003444445455555565666777777777888888889899999999A9AAAAAAAAAABB73234323232222222222222222222222002220200022222202002000202222202000000000000200000022220200000000000000000000202002020002200000000222200020200002000000000000000200220022000000000000002000000200000020002002000020000000000000202000000200000000222202020023320000022022222002000020022020222000000000000202020222222202222222223237CCCCCCCBCCBCCCBCCCCCBCBCCCCCCBCCBCCBCCBBBBBAA99887755543322020000000000000000000000000000000000000;
		rom_data[373] <= 3840'h55555556666777777778888888888999999A9A9AAAAAAAAAAABC8423322222232223222222222222222222002002020223320202002022222200200202000000002000220202202000200000200000000000020002200000000000020000000000000200200000000002000000000000000000000000002000020000000022000000020000002200000002002000002220000022200020002222000202020020222000220000020222200000200000202020202332222222222222325ACCCCBCCCCCCCBBCBCBCBCCCCCCBCBCCBCBCCCBCBBBA99887765553332202000000000000000000000000000000000000004444445555555556666777777778888888888999999A9A9AAAAAAAAAAABC8423322222232223222222222222222222002002020223320202002022222200200202000000002000220202202000200000200000000000020002200000000000020000000000000200200000000002000000000000000000000000002000020000000022000000020000002200000002002000002220000022200020002222000202020020222000220000020222200000200000202020202332222222222222325ACCCCBCCCCCCCBBCBCBCBCCCCCCBCBCCBCBCCCBCBBBA9988776555333220200000000000000000000000000000000000000;
		rom_data[374] <= 3840'h55555565666777777778888888889889999999999AAAAAAAAABB9532232323222222222332222222332220000200200223322202202020202022020020200000000020220023220000002000002000000000000000020002000022000000000000220000200002000200022000000000000000000000000000000000000000002020000000000020000020000000000220000222202202000200200020222202202202000020202022000000002002022202022332222220222003437CCCBCCBCCBCBCCCCBCBCCCCCBCCCBCCBCBCBBBBBBBAA99877655433220200000000000000000000000000000000000000004344545455555565666777777778888888889889999999999AAAAAAAAABB9532232323222222222332222222332220000200200223322202202020202022020020200000000020220023220000002000002000000000000000020002000022000000000000220000200002000200022000000000000000000000000000000000000000002020000000000020000020000000000220000222202202000200200020222202202202000020202022000000002002022202022332222220222003437CCCBCCBCCBCBCCCCBCBCCCCCBCCCBCCBCBCBBBBBBBAA9987765543322020000000000000000000000000000000000000000;
		rom_data[375] <= 3840'h55555555666677777788888888888999999A9A9AAAAAAAAAAABBA733232333222332222230222222332020200200020222432022222020202202222202000000002002200223220020020000000200000000000000000020000000002200000000020200000020000000000000200000000000000000000000002000000002000020000000000020200000202020000200020022022320200202002222202022022002220202202000202220000000202020222222222222220024459CCCCCCCCBCCCCBCBCCCCCCCBCCBCBCBCBCBCCBBBAA9988775544332200000000000000000000020000000000000000000003444445555555555666677777788888888888999999A9A9AAAAAAAAAAABBA733232333222332222230222222332020200200020222432022222020202202222202000000002002200223220020020000000200000000000000000020000000002200000000020200000020000000000000200000000000000000000000002000000002000020000000000020200000202020000200020022022320200202002222202022022002220202202000202220000000202020222222222222220024459CCCCCCCCBCCCCBCBCCCCCCCBCCBCBCBCBCBCCBBBAA998877554433220000000000000000000002000000000000000000000;
		rom_data[376] <= 3840'h55555565666677777778888888888899999999A9AAAAAAAAAAAAB84323323232233222222202222023220020020020202352200002200002222020000020000000000000000202200000000000000002000000000000020002202000000200000000000000000000000000000000000000202000000000002000000002200200200000000200000020220020020020002002022220542000002000022020020222022020002020020002430000000200022022202222322220202547BCCBCBCBCCCCBCCCCCBBCCBCCCCCCCBCCCBCCBBBAA99887765443222020000000000000000002202200000000000000000003444444555555565666677777778888888888899999999A9AAAAAAAAAAAAB84323323232233222222202222023220020020020202352200002200002222020000020000000000000000202200000000000000002000000000000020002202000000200000000000000000000000000000000000000202000000000002000000002200200200000000200000020220020020020002002022220542000002000022020020222022020002020020002430000000200022022202222322220202547BCCBCBCBCCCCBCCCCCBBCCBCCCCCCCBCCCBCCBBBAA9988776544322202000000000000000000220220000000000000000000;
		rom_data[377] <= 3840'h5555555566677777788888888888999999999A9AAAAAAAAAAAABB95233232223222222222222220222222020000202202222202020000023300020002220000000000002002202000000002000000000200000000000200000002000002000000000002000000200000000000000002020002000000000202220000022200000000000000000020000000002000002000020022222432002020200220200022022220200022020200000200002002020202020202222222222023549CCCCCCCCCBCCCCBCBCCCCBCCBCBCBCBCBCCBBBAAA99887755443220000000000000000000022222202000000000000000000444445455555555566677777788888888888999999999A9AAAAAAAAAAAABB95233232223222222222222220222222020000202202222202020000023300020002220000000000002002202000000002000000000200000000000200000002000002000000000002000000200000000000000002020002000000000202220000022200000000000000000020000000002000002000020022222432002020200220200022022220200022020200000200002002020202020202222222222023549CCCCCCCCCBCCCCBCBCCCCBCCBCBCBCBCBCCBBBAAA99887755443220000000000000000000022222202000000000000000000;
		rom_data[378] <= 3840'h5555556566767777777888888889888999999999AAAAAAAAAABABA733232222222222222222222220222220202000222022220002222002332220200022000000000000000020000000200222000002000000000000000000002000000000200000020000000000000000000000000220000000000000000222000000000000002000002000020000200000222000002000022222222020020000202020200222202200000000002000002000000200220202202022222222202436BCBCBBCCBCCCCBCCBCBCBCCBCCCCCCBCBCBCBBBAA998877555332202000000000000000000222332322200000000000000000344444555555556566767777777888888889888999999999AAAAAAAAAABABA733232222222222222222222220222220202000222022220002222002332220200022000000000000000020000000200222000002000000000000000000002000000000200000020000000000000000000000000220000000000000000222000000000000002000002000020000200000222000002000022222222020020000202020200222202200000000002000002000000200220202202022222222202436BCBCBBCCBCCCCBCCBCBCBCCBCCCCCCBCBCBCBBBAA998877555332202000000000000000000222332322200000000000000000;
		rom_data[379] <= 3840'h555555566667777778788888888889989999A9A9AAAAAAAAAAAABB953232322222222222222022222202020000200200200202020022000022220200000000000000000222200002202000200000200000000000200000002020200000000000000000000000000000002000000002000000000000000000000200000200000000000000000000000000000232200000000222202000000202000202020233322022000000000000000200000002022020202020222220232022449CCCCCCCCCCBCCCCBCCBCCBCCCCBCBBCCCBCBBBAA998877554332200000000000000000002233434333220000000000000000044444555555555566667777778788888888889989999A9A9AAAAAAAAAAAABB953232322222222222222022222202020000200200200202020022000022220200000000000000000222200002202000200000200000000000200000002020200000000000000000000000000000002000000002000000000000000000000200000200000000000000000000000000000232200000000222202000000202000202020233322022000000000000000200000002022020202020222220232022449CCCCCCCCCCBCCCCBCCBCCBCCCCBCBBCCCBCBBBAA9988775543322000000000000000000022334343332200000000000000000;
		rom_data[380] <= 3840'h55555556666777777788888888898989999999A9AAAAAAAAAAAAABA6333332232220222022220222222222020022002000202002000000000022200000000000000000002002002020000000000000000000000000000000002200000000000000000000002000000000000000000200000000000000000002000002020002000000000000000000000000022220200000002020000000002020020202223322220200020020000000000000000000002022200223202222202247CCBCBCCBCBCCCBCBCCCCBCCCBCCCBCBCBCCBBBA9988876554332220000000000000000022334455544333200000000000000004444444555555556666777777788888888898989999999A9AAAAAAAAAAAAABA6333332232220222022220222222222020022002000202002000000000022200000000000000000002002002020000000000000000000000000000000002200000000000000000000002000000000000000000200000000000000000002000002020002000000000000000000000000022220200000002020000000002020020202223322220200020020000000000000000000002022200223202222202247CCBCBCCBCBCCCBCBCCCCBCCCBCCCBCBCBCCBBBA998887655433222000000000000000002233445554433320000000000000000;
		rom_data[381] <= 3840'h555555665667777778888888888889899999A99AAAAAAAAAAAABABB843233222222222222220220223202200022220002002020000020000020202200000000000000000000220002000220202000000000000000000000000200000000020000000000000000000000000000000000000000000000000000000002000020200000000000000000000000000020200000002220020000000202022202002222232002000000000000000000000000202020020222222220002236BCCCCCCBCCCCBCCBCBCBCCCBBCCCBCBCCCCBBAA998877755433220000000000000000022334555655555433200000000000000043444555555555665667777778888888888889899999A99AAAAAAAAAAAABABB843233222222222222220220223202200022220002002020000020000020202200000000000000000000220002000220202000000000000000000000000200000000020000000000000000000000000000000000000000000000000000000002000020200000000000000000000000000020200000002220020000000202022202002222232002000000000000000000000000202020020222222220002236BCCCCCCBCCCCBCCBCBCBCCCBBCCCBCBCCCCBBAA9988777554332200000000000000000223345556555554332000000000000000;
		rom_data[382] <= 3840'h5555555666677777787888888889889999999A99A9AAAAAAAAAABBB953333322332022232022202223222220202222000202020200000200022020220000000000000000220020000200020000000000000000000000000000000200000000000000020000000000000000020000000000000000200000000000000000022200000000200000000000000000000000000002222000000020000202020202020220200200000002000000000000000022002020222222222002249CCCBCBCCCCBCCCCCCCCCCCBCCCCBCBCBBCBBBA99887765543222200000000000000022234455777777655432000000000000000444544555555555666677777787888888889889999999A99A9AAAAAAAAAABBB953333322332022232022202223222220202222000202020200000200022020220000000000000000220020000200020000000000000000000000000000000200000000000000020000000000000000020000000000000000200000000000000000022200000000200000000000000000000000000002222000000020000202020202020220200200000002000000000000000022002020222222222002249CCCBCBCCCCBCCCCCCCCCCCBCCCCBCBCBBCBBBA99887765543222200000000000000022234455777777655432000000000000000;
		rom_data[383] <= 3840'h5555556566677777788888888888998999999A9A9AAAAAAAAAABABBA7333322222222233320222022222220200022002020222200000200000020200020000000000000020020000202000000000000002000000000000000000000000000000000000000000000000000002000000000000000000000000000000000002320000000000000000000000000000000000020222022020000020002000002020020200000200202000002000000002020002002022220220022225ACCCCCCCBCCCCBCBCBCBCCBCCBBCCCCBBCBBAAA98776554432220000000000000000223445567788888776543200000000000000344445555555556566677777788888888888998999999A9A9AAAAAAAAAABABBA7333322222222233320222022222220200022002020222200000200000020200020000000000000020020000202000000000000002000000000000000000000000000000000000000000000000000002000000000000000000000000000000000002320000000000000000000000000000000000020222022020000020002000002020020200000200202000002000000002020002002022220220022225ACCCCCCCBCCCCBCBCBCBCCBCCBBCCCCBBCBBAAA98776554432220000000000000000223445567788888776543200000000000000;
		rom_data[384] <= 3840'h5555555666677777777888888888989899999A99A9AAAAAAAAAABABB9533333222222223222222222222222202000202002202022000020020002022000000000000000000000000220200000000000000000000000000002000000200000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000222002000202002220000002002020020002000000000000200000020020200202202202222002225ACCBCCBCCCCBCCCCCCCCBCCCBCCCBCBCBBBBA9988766544322202000000000000022334556778899999887543200000000000000444444455555555666677777777888888888989899999A99A9AAAAAAAAAABABB9533333222222223222222222222222202000202002202022000020020002022000000000000000000000000220200000000000000000000000000002000000200000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000222002000202002220000002002020020002000000000000200000020020200202202202222002225ACCBCCBCCCCBCCCCCCCCBCCCBCCCBCBCBBBBA9988766544322202000000000000022334556778899999887543200000000000000;
		rom_data[385] <= 3840'h5555555566677777788888888888898999999A9A9AAAAAAAAAAAAABBA833223222222022222020222202223220020020022022020020200200022000000000000000000020200020000000000000000002200000000200000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000002200000000000000000000002222000000020202000002002020002000202000200000020000200200002020222022020200222235BCCCCBCCBCCCCBCCCBCCCCBCCBCBCBCBBBBAA988765544322200000000000000022345557788999AABA987653320000000000000444454555555555566677777788888888888898999999A9A9AAAAAAAAAAAAABBA833223222222022222020222202223220020020022022020020200200022000000000000000000020200020000000000000000002200000000200000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000002200000000000000000000002222000000020202000002002020002000202000200000020000200200002020222022020200222235BCCCCBCCBCCCCBCCCBCCCCBCCBCBCBCBBBBAA988765544322200000000000000022345557788999AABA987653320000000000000;
		rom_data[386] <= 3840'h5555555666677777778888888888989899999999A9AAAAAAAAAAABABBA52233222202222220202222222222220000200000020202000220000000220000000000000000000202020222000000000000000200000020022000000000000000000000000000000000000000000000000000000000000000000000002000002200000000000002000000000000000000000000220200000203322020200022020020000000000020000020020000000200000222002222220222335BCCBCCCCCCCBCCBCBCBCBBCBCCBCCCCBBAA9998775544222200000000000000023344567788999AABBBA88654320000000000000444454555555555666677777778888888888989899999999A9AAAAAAAAAAABABBA52233222202222220202222222222220000200000020202000220000000220000000000000000000202020222000000000000000200000020022000000000000000000000000000000000000000000000000000000000000000000000002000002200000000000002000000000000000000000000220200000203322020200022020020000000000020000020020000000200000222002222220222335BCCBCCCCCCCBCCBCBCBCBBCBCCBCCCCBBAA9998775544222200000000000000023344567788999AABBBA88654320000000000000;
		rom_data[387] <= 3840'h5555555666677777778888888888898999999A9A9AAAAAAAAAAABAABBB73233322222222222202220222222220000002020222200220200000002200000000000000000002202000200200000000000000000000000020200000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000002202000002023220000002020220000200000200000000200200000002002020200222222202233336BCCCCBCBCCCCBCCCCCCBCCBCBCCCBBBBAA99987755433220000000000000000233455777889AAABBBBBA98754320000000000000344445455555555666677777778888888888898999999A9A9AAAAAAAAAAABAABBB73233322222222222202220222222220000002020222200220200000002200000000000000000002202000200200000000000000000000000020200000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000002202000002023220000002020220000200000200000000200200000002002020200222222202233336BCCCCBCBCCCCBCCCCCCBCCBCBCCCBBBBAA99987755433220000000000000000233455777889AAABBBBBA98754320000000000000;
		rom_data[388] <= 3840'h5555555666767777777888888888889899999999A9AAAAAAAAAAAAAABB94323322222222222202022022222222200000002020222020020000000200000000000000000000020200200200000000000000000000000000000000000000000000000000000000000000220000000000000000000000000000000000002000000000000000000000000000000000000000002020020000222020020200000000020000000000000000020000000000020202220202022222233335CCBBCCCCCCBCCBCBBCBCBBCBCCBBBBBAA9988765543320200000000000000223445677889AAABBBBBBBA98765330000000000000444444555555555666767777777888888888889899999999A9AAAAAAAAAAAAAABB94323322222222222202022022222222200000002020222020020000000200000000000000000000020200200200000000000000000000000000000000000000000000000000000000000000220000000000000000000000000000000000002000000000000000000000000000000000000000002020020000222020020200000000020000000000000000020000000000020202220202022222233335CCBBCCCCCCBCCBCBBCBCBBCBCCBBBBBAA9988765543320200000000000000223445677889AAABBBBBBBA98765330000000000000;
		rom_data[389] <= 3840'h555555565666777777788888888889989999A99A9AAAAAAAAAAAAAAABBA7322222222222222202020222022202000000202020220200000000020000000000000000000000002002000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000002002000020000000000000000000000000000000000000000200200022020200200000200000000202000020000000000000000020002020022222022223333235CCCCBCCCBCCCBCCBCBCBCCCCBCBBBBAA9988765543322000000000000000233445678899AABBBBBBBBBAA876542200000000000044444555555555565666777777788888888889989999A99A9AAAAAAAAAAAAAAABBA7322222222222222202020222022202000000202020220200000000020000000000000000000000002002000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000002002000020000000000000000000000000000000000000000200200022020200200000200000000202000020000000000000000020002020022222022223333235CCCCBCCCBCCCBCCBCBCBCCCCBCBBBBAA9988765543322000000000000000233445678899AABBBBBBBBBAA8765422000000000000;
		rom_data[390] <= 3840'h5555555566667777777788888888898999999A9AAAAAAAAAAAAAAAABABB9522323222222232220202202202222020000020002002020000000002000000000000000000020200000200200000000000000000000000000000200000000000000000200000000000000033200000000000000000000000000000000200200000000000000000000000000000000000000002000000000200000020000022000020000000000200000002000000000200022022022202233433336CCCCCCBCCBCBCCBCCCCCCBCBCCBBBAA9887765443222000000000000002233455678899ABBBBBBBBBBBAA8775430000000000000444454455555555566667777777788888888898999999A9AAAAAAAAAAAAAAAABABB9522323222222232220202202202222020000020002002020000000002000000000000000000020200000200200000000000000000000000000000200000000000000000200000000000000033200000000000000000000000000000000200200000000000000000000000000000000000000002000000000200000020000022000020000000000200000002000000000200022022022202233433336CCCCCCBCCBCBCCBCCCCCCBCBCCBBBAA9887765443222000000000000002233455678899ABBBBBBBBBBBAA8775430000000000000;
		rom_data[391] <= 3840'h5555555666667777777888888888899999999A9AAAAAAAAAAAAAAABAABBB732232322220223202202020222022200200000022020220200200000000000000000000000000002020002020220000000000000000000000000020000000000000000200000000000000022200000000000000000000000000000000000000000000000000000000000000000020000000002000002220002020200002200020000202000202000000002000020000002022220222222233443337CBCBCCCCCCBCBCCBCBBBBCBCBBBBAA988776544322000000000000000223345577889ABBBBCBBBBBBBBAA9875422000000000000344444555555555666667777777888888888899999999A9AAAAAAAAAAAAAAABAABBB732232322220223202202020222022200200000022020220200200000000000000000000000000002020002020220000000000000000000000000020000000000000000200000000000000022200000000000000000000000000000000000000000000000000000000000000000020000000002000002220002020200002200020000202000202000000002000020000002022220222222233443337CBCBCCCCCCBCBCCBCBBBBCBCBBBBAA988776544322000000000000000223345577889ABBBBCBBBBBBBBAA9875422000000000000;
		rom_data[392] <= 3840'h55555555666667777777888888889899999999AAAAAAAAAAAAAAAAABABBC852232322222222222222202022222220000000002002002200000000200000000000000000000000022002022200000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000202020000200000000000000000000000000000000000202200020200202202000000220200020220200200000000002202002200200202022222223343344337CCCCCCCBCBCCCCBCBCCCCBBBBBAA9988775544322200000000000000233455678899AABBBBBBBBBBBBBB998754300000000000004444454555555555666667777777888888889899999999AAAAAAAAAAAAAAAAABABBC852232322222222222222202022222220000000002002002200000000200000000000000000000000022002022200000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000202020000200000000000000000000000000000000000202200020200202202000000220200020220200200000000002202002200200202022222223343344337CCCCCCCBCBCCCCBCBCCCCBBBBBAA9988775544322200000000000000233455678899AABBBBBBBBBBBBBB99875430000000000000;
		rom_data[393] <= 3840'h5555555666667777777888888888899999999A9AAAAAAAAAAAAAABABABABB73223222222222022320222022020202020000000020220000000000000020000000000000000200000000000000000000000000000000002200000000000000000000000000002000000000000000000000000000000000000000000200000000200000000000000000000000022000000020000200200023300022020000000002300020000000000000002020000020222222202234444443237CCBCBCCCCCBCBCCCCBCBBBBBBAA9988775543322000000000000002233455678899AABBBBBBBBBBBBBBAA8875432000000000000444445455555555666667777777888888888899999999A9AAAAAAAAAAAAAABABABABB73223222222222022320222022020202020000000020220000000000000020000000000000000200000000000000000000000000000000002200000000000000000000000000002000000000000000000000000000000000000000000200000000200000000000000000000000022000000020000200200023300022020000000002300020000000000000002020000020222222202234444443237CCBCBCCCCCBCBCCCCBCBBBBBBAA9988775543322000000000000002233455678899AABBBBBBBBBBBBBBAA8875432000000000000;
		rom_data[394] <= 3840'h5555555566667777777888888888898999999A99AAAAAAAAAAAAAAAAAABAC85223322220222202222020202220200200000002000022000000000002000000000000000002002020000002000000000000000000000000200000000000000000000000000020000000000000000000000000000000000000000020000000000000000000000000000000000003300000020020202002022222000000020202002202000200000000002000002000002000223220355544432227CCCCCCBCBCCBCBBBCBCBCBBBAA9988765543322200000000000002234456778899ABBBBBBBBBBBBBBBBBA9875542000000000000444445455555555566667777777888888888898999999A99AAAAAAAAAAAAAAAAAABAC85223322220222202222020202220200200000002000022000000000002000000000000000002002020000002000000000000000000000000200000000000000000000000000020000000000000000000000000000000000000000020000000000000000000000000000000000003300000020020202002022222000000020202002202000200000000002000002000002000223220355544432227CCCCCCBCBCCBCBBBCBCBCBBBAA9988765543322200000000000002234456778899ABBBBBBBBBBBBBBBBBA9875542000000000000;
		rom_data[395] <= 3840'h55555565666677777787888888889899999999A9AAAAAAAAAAAAAAABABABBB7322232220222222220222022220002002000000220002000000000020022000000000000000020000000200200000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000020000000000000000000000000000020000222200000000200202000202000000020200022002020000000000000000000200002222220222202466454322037CCCCCCCBCCCCCCCBCBCBBBBBA998876554332200000000000000333455677889AAABBBBBBCBBCBBBBBBBA98765432000000000004445445555555565666677777787888888889899999999A9AAAAAAAAAAAAAAABABABBB7322232220222222220222022220002002000000220002000000000020022000000000000000020000000200200000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000020000000000000000000000000000020000222200000000200202000202000000020200022002020000000000000000000200002222220222202466454322037CCCCCCCBCCCCCCCBCBCBBBBBA998876554332200000000000000333455677889AAABBBBBBCBBCBBBBBBBA9876543200000000000;
		rom_data[396] <= 3840'h555555556666777777888888888888999999A9A9AAAAAAAAAAAAAAAAAABABC9423222222222202202222202220220002000000000000200000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000020000000000000000000000000000000000020002020000000200020000202002000202000000000000000200020200232002222022455554222038CCCCCCBCBCBCCBCBCBCBBBBAA98876544322200000000000002233455778899AABCBBBBBBBBBBBBBBBBBA988755332220000000044444454555555556666777777888888888888999999A9A9AAAAAAAAAAAAAAAAAABABC9423222222222202202222202220220002000000000000200000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000020000000000000000000000000000000000020002020000000200020000202002000202000000000000000200020200232002222022455554222038CCCCCCBCBCBCCBCBCBCBBBBAA98876544322200000000000002233455778899AABCBBBBBBBBBBBBBBBBBA9887553322200000000;
		rom_data[397] <= 3840'h555555556666777777888888888899899999999AAAAAAAAAAAAAABABAAABBBA732223222020222202020202220200202000000022020000000000002000220000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000200200200200020002222000000000000000000000000000000000220202220202202224545542222048EBCBCCCCCCCBCBCCBCBBBBAA98776554322000000000000002234555788899AABBBBBBBBBBBBBBBBBBBBBA98775543323232220244445454555555556666777777888888888899899999999AAAAAAAAAAAAAABABAAABBBA732223222020222202020202220200202000000022020000000000002000220000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000200200200200020002222000000000000000000000000000000000220202220202202224545542222048EBCBCCCCCCCBCBCCBCBBBBAA98776554322000000000000002234555788899AABBBBBBBBBBBBBBBBBBBBBA987755433232322202;
		rom_data[398] <= 3840'h55555555566677777778888888888899999A99A9AAAAAAAAAAAAAAAAABABABB84232222222222222202020002022000022000000022220000000000000022000000000000000000000000000000000000000000000000000000002200000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000202000200200200222000200200000000000000000000000000200202020202020224554442222224ACCCCCCCCBCBCCCCBCBCBAA99887655432200000000000000234455678889AAABBBBCBBBCBBBBBBCBBBBBAA9987755544443333334444454555555555566677777778888888888899999A99A9AAAAAAAAAAAAAAAAABABABB84232222222222222202020002022000022000000022220000000000000022000000000000000000000000000000000000000000000000000000002200000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000202000200200200222000200200000000000000000000000000200202020202020224554442222224ACCCCCCCCBCBCCCCBCBCBAA99887655432200000000000000234455678889AAABBBBCBBBCBBBBBBCBBBBBAA998775554444333333;
		rom_data[399] <= 3840'h555555556566777778888888888899899999999AAAAAAAAAAAAAAAAAAAAAABBA7423222220222022020202202020022020200000223200020000000000000200000000000000000000000000000000000000000000000000000002222000000000000000000000000000000020000000000000000000000200000000000000000000000000000000000000000000000202000002022000000000002000000000000020000000000000000020000202020202235554422020025CCCBCBCBCCBCBBBCBCBBBA99887754432200000000000000233455678899AABBBBBBBBBBBBBCBBBBBBBBBBBA9888776555554444444444555555555556566777778888888888899899999999AAAAAAAAAAAAAAAAAAAAAABBA7423222220222022020202202020022020200000223200020000000000000200000000000000000000000000000000000000000000000000000002222000000000000000000000000000000020000000000000000000000200000000000000000000000000000000000000000000000202000002022000000000002000000000000020000000000000000020000202020202235554422020025CCCBCBCBCCBCBBBCBCBBBA99887754432200000000000000233455678899AABBBBBBBBBBBBBCBBBBBBBBBBBA98887765555544444;
		rom_data[400] <= 3840'h555555556666777777888888888888999999A9A9AAAAAAAAAAAAAABABAABBBBB9632322222202222202020202202022220200000022020002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000222000000000000000000002200000022000000002000000000000000000000000000000200200200200200000000000020000000000000000000000000000002002020220222355555322022027ECCCCCCCCCCCCCBBBBBAA9988765543220000000000000223445577889AABBBBBBCBBBBBBBBBBBBBBBBBBBBAA998877767766565544445455555555556666777777888888888888999999A9A9AAAAAAAAAAAAAABABAABBBBB9632322222202222202020202202022220200000022020002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000222000000000000000000002200000022000000002000000000000000000000000000000200200200200200000000000020000000000000000000000000000002002020220222355555322022027ECCCCCCCCCCCCCBBBBBAA9988765543220000000000000223445577889AABBBBBBCBBBBBBBBBBBBBBBBBBBBAA9988777677665655;
		rom_data[401] <= 3840'h55555556666677777888888888899999999A99A9AAAAAAAAAAAAAAABAABABABBB83333222022222322022222022022332020000002000000000000000000000000000000000000020000000000000000000000000000000000000000000020000000000000000000000000022000000000000000000000220000002200000000000000000000000000000000000000200000000000200000000002000000000000000000000000020000002002022222222345555432222004ACCCCCCCCBCBBBCCBBBAA9987765543220000000000000033355678889AABBBBBCBBBBBCBBBBBBBBBCBBBBBBAAA9988888887777774444545555555556666677777888888888899999999A99A9AAAAAAAAAAAAAAABAABABABBB83333222022222322022222022022332020000002000000000000000000000000000000000000020000000000000000000000000000000000000000000020000000000000000000000000022000000000000000000000220000002200000000000000000000000000000000000000200000000000200000000002000000000000000000000000020000002002022222222345555432222004ACCCCCCCCBCBBBCCBBBAA9987765543220000000000000033355678889AABBBBBCBBBBBCBBBBBBBBBCBBBBBBAAA998888888777777;
		rom_data[402] <= 3840'h555555556666777777788888888889899999A9A9AAAAAAAAAAAAAAAAABABBBBBBA5223222222022202000222020202222200000000022002000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000200020000000022200000000000000020000000200002000020202200222455654322222026ECCCCCCBCCCCCCBBBBAA9988775533220000000000000223455678899ABBBBCBBBBBBBBBBCBBBBBBBBBBBBBBBAAAA999998988888844454555555555556666777777788888888889899999A9A9AAAAAAAAAAAAAAAAABABBBBBBA5223222222022202000222020202222200000000022002000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000200020000000022200000000000000020000000200002000020202200222455654322222026ECCCCCCBCCCCCCBBBBAA9988775533220000000000000223455678899ABBBBCBBBBBBBBBBCBBBBBBBBBBBBBBBAAAA9999989888888;
		rom_data[403] <= 3840'h555555566667777777788888888898999999999AAAAAAAAAAAAAAAAAAABBABABBB742332222222020202022202022002002200000002002002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000200000000000000000000000000000000000000020000000022020200200200000000002200000000000000000000000200000002020022002233556665432222005ACCCCCCCCCBCCBBCBBAA9988765543322000000000000223445678889AABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABAAAAAAA9A99989944454555555555566667777777788888888898999999999AAAAAAAAAAAAAAAAAAABBABABBB742332222222020202022202022002002200000002002002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000200000000000000000000000000000000000000020000000022020200200200000000002200000000000000000000000200000002020022002233556665432222005ACCCCCCCCCBCCBBCBBAA9988765543322000000000000223445678889AABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABAAAAAAA9A999899;
		rom_data[404] <= 3840'h555555556667777777888888888989999999A9A9AAAAAAAAAAAAAAAABAAABABABBA63222222222202022200220200200220000000000200000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002200000000000000000000000000000000000000000000000000222000020000000000000000002020000000000000000000000000000000200202222235787665322220239ECCCCCCCCCCCBCBBBAA9988765543222000000000000233445778899ABBBBBBBBBBBBBBBBBBBBCBBCBBBBBBBBBBBBBBBBAABAAAAA9A44545555555555556667777777888888888989999999A9A9AAAAAAAAAAAAAAAABAAABABABBA63222222222202022200220200200220000000000200000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002200000000000000000000000000000000000000000000000000222000020000000000000000002020000000000000000000000000000000200202222235787665322220239ECCCCCCCCCCCBCBBBAA9988765543222000000000000233445778899ABBBBBBBBBBBBBBBBBBBBCBBCBBBBBBBBBBBBBBBBAABAAAAA9A;
		rom_data[405] <= 3840'h55555556666777777788888888888999999A9A9AAAAAAAAAAAAAAAAAAAABABAABBB94222222222022220200002020222202200000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000002000000000000000000000000000000000000000000000000000000000200200000020200000000000000000000200000000000000000020202202022246CB875532322249CCCCCCCCCCCCBCBBBA99887765543320000000000000223445678899ABBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBABA4445545555555556666777777788888888888999999A9A9AAAAAAAAAAAAAAAAAAAABABAABBB94222222222022220200002020222202200000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000002000000000000000000000000000000000000000000000000000000000200200000020200000000000000000000200000000000000000020202202022246CB875532322249CCCCCCCCCCCCBCBBBA99887765543320000000000000223445678899ABBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBABA;
		rom_data[406] <= 3840'h555555566666777778788888888889899999A9A9AAAAAAAAAAAAAABABAAAAAABABBB7322222222202020200200200000000220000000020020200000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000200000002300000000200000000000000000002000200000020002022222335998754222235ACCCCCCCCCCCCCBBBBAA9987765443222000000000000233455778899ABBBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB44545555555555566666777778788888888889899999A9A9AAAAAAAAAAAAAABABAAAAAABABBB7322222222202020200200200000000220000000020020200000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000200000002300000000200000000000000000002000200000020002022222335998754222235ACCCCCCCCCCCCCBBBBAA9987765443222000000000000233455778899ABBBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[407] <= 3840'h55555566667777777788888888899899999A9A9AAAAAAAAAAAAAAAAABABBBBBABBBB952222323322020200202002020200220200000000002000000002000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000200000002000000000000200000000000000002202020020202233434887543458BCCCCCCCCCCCCBCBBBA9988776544322000000000000023345677889AABBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB4545555555555566667777777788888888899899999A9A9AAAAAAAAAAAAAAAAABABBBBBABBBB952222323322020200202002020200220200000000002000000002000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000200000002000000000000200000000000000002202020020202233434887543458BCCCCCCCCCCCCBCBBBA9988776544322000000000000023345677889AABBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[408] <= 3840'h55555566676777777788888888888989999999A9AAAAAAAAAAAAAAAAAAAAAAABBAABB852222233202020220202002002200020000000000002000000022000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000002000000000000000000020000000000202022222022232259CA989ABECCCCCCCCCCCCCCBBAAA988776544322200000000000223445577899AAABBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB4455555555555566676777777788888888888989999999A9AAAAAAAAAAAAAAAAAAAAAAABBAABB852222233202020220202002002200020000000000002000000022000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000002000000000000000000020000000000202022222022232259CA989ABECCCCCCCCCCCCCCBBAAA988776544322200000000000223445577899AAABBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[409] <= 3840'h555555656677777777788888888998999999A99AAAAAAAAAAAAAAAAAAAABABABAABABB7322222222022202020002220220020200000000002020000000200000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200020000000000000000000000000000000000002020002020202220020222038CCCECECCCCCCCCCCCCCCCBBBAA9988775543322000000000000023345578889AABBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB55455555555555656677777777788888888998999999A99AAAAAAAAAAAAAAAAAAAABABABAABABB7322222222022202020002220220020200000000002020000000200000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200020000000000000000000000000000000000002020002020202220020222038CCCECECCCCCCCCCCCCCCCBBBAA9988775543322000000000000023345578889AABBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[410] <= 3840'h5555556667677777777888888898899999A999A9AAAAAAAAAAAAAAAAAAAAAABBBABABB952232222222022202020022000200020000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200200000000000000000000000000000000000200000000200020202022027CCCCCCCCCCCCCCCCCCCBBCBBAA9988765543322200000000000223355677889AABBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB445555555555556667677777777888888898899999A999A9AAAAAAAAAAAAAAAAAAAAAABBBABABB952232222222022202020022000200020000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200200000000000000000000000000000000000200000000200020202022027CCCCCCCCCCCCCCCCCCCBBCBBAA9988765543322200000000000223355677889AABBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[411] <= 3840'h5555556666767777778888888888999999999A9AAAAAAAAAAAAAAAAAAABBBABBBABAABB8423222202022200200202022202000020000000000020000002000000000000000000000000000000000000000000000000000022000000000000000000000000030000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000002000202002220020024BCCCCCCCCCCCCCCCCBCBCCBBBA9988765543320000000000000223345678899ABBBBBBBBBBBBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB545555555555556666767777778888888888999999999A9AAAAAAAAAAAAAAAAAAABBBABBBABAABB8423222202022200200202022202000020000000000020000002000000000000000000000000000000000000000000000000000022000000000000000000000000030000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000002000202002220020024BCCCCCCCCCCCCCCCCBCBCCBBBA9988765543320000000000000223345678899ABBBBBBBBBBBBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[412] <= 3840'h555556666677777778888888888889899999A999AAAAAAAAAAAAAAAAAAAAABAAABABABBA732222222020220022000202020000000000000020002000000200000000000000000000000000000000000000000000000000022000000000000000000000000200000000000000000000220000000000000000000000000000000000000000000000000000000000000000200000000000000000200020000000000000000000020000200202000222002239CCCCCCCCCCCCCCCCCCBCBCBBA9988775543222200000000000223455677889AABBBBBBBCBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB45555555555556666677777778888888888889899999A999AAAAAAAAAAAAAAAAAAAAABAAABABABBA732222222020220022000202020000000000000020002000000200000000000000000000000000000000000000000000000000022000000000000000000000000200000000000000000000220000000000000000000000000000000000000000000000000000000000000000200000000000000000200020000000000000000000020000200202000222002239CCCCCCCCCCCCCCCCCCBCBCBBA9988775543222200000000000223455677889AABBBBBBBCBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[413] <= 3840'h5556666667777777788888888888899999999A9AAAAAAAAAAAAAAAAAAAAAAAABAAAAAABB95322220202020202020200200020200200000020202000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000020200200022220202038CCCCCCCCCCCCCCCCCCBCBBBBAA988775543322000000000000023345677899ABBBBBBCBBBCBBBBBBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB455555555556666667777777788888888888899999999A9AAAAAAAAAAAAAAAAAAAAAAAABAAAAAABB95322220202020202020200200020200200000020202000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000020200200022220202038CCCCCCCCCCCCCCCCCCBCBBBBAA988775543322000000000000023345677899ABBBBBBCBBBCBBBBBBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[414] <= 3840'h55556566667777777788888888888989999999A9AAAAAAAAAAAAAAAAAAABABBABABABABBB842222220200202000002002020022000002000002002000000002002000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000200200000202025AECCBCCCCCCCCCCCCCCCCBBBAA988765543220000000000000223455678899AABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB5555555555556566667777777788888888888989999999A9AAAAAAAAAAAAAAAAAAABABBABABABABBB842222220200202000002002020022000002000002002000000002002000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000200200000202025AECCBCCCCCCCCCCCCCCCCBBBAA988765543220000000000000223455678899AABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[415] <= 3840'h5556666666777777788888888888899999999A9AAAAAAAAAAAAAAAAAABABAAAAABABABABBA73222220202000020220002000202220202000000020000000020000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002200000020000000000000000000000000000000000000000000000000000000000020002020202020227BCCCCCCCCCCCCCCCCCCBCBBAA988775543320000000000000223445678899ABBBBBBBCBBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB545555555556666666777777788888888888899999999A9AAAAAAAAAAAAAAAAAABABAAAAABABABABBA73222220202000020220002000202220202000000020000000020000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002200000020000000000000000000000000000000000000000000000000000000000020002020202020227BCCCCCCCCCCCCCCCCCCBCBBAA988775543320000000000000223445678899ABBBBBBBCBBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[416] <= 3840'h55556566777677778788888888898999999999A9AAAAAAAAAAAAAAAAAAAAAAABAAAABAAAABA5322222202022200020200220002220020200000002000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000022200002200000000000000000200002000000002000000000000000000000020000002200020020202236ACCCCCCBCCCCCCCBBCCBBBAA998775543220200000000000223445677899ABBBBBBBBBCBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB5555555555556566777677778788888888898999999999A9AAAAAAAAAAAAAAAAAAAAAAABAAAABAAAABA5322222202022200020200220002220020200000002000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000022200002200000000000000000200002000000002000000000000000000000020000002200020020202236ACCCCCCBCCCCCCCBBCCBBBAA998775543220200000000000223445677899ABBBBBBBBBCBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[417] <= 3840'h566666666767777778888888888899999999A9A9AAAAAAAAAAAAAAAAAABAAAAAABABAAAAABB8422202220202200020002000000202000000000000000000002000020000000000000000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000000000000000000000000000000000002200000000000000002200022000000020020000000000000000000000200022200200200222236BCCCCCCCCBCCCCCCCCBBBAA988775543322000000000000223445678889AABBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB55555555566666666767777778888888888899999999A9A9AAAAAAAAAAAAAAAAAABAAAAAABABAAAAABB8422202220202200020002000000202000000000000000000002000020000000000000000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000000000000000000000000000000000002200000000000000002200022000000020020000000000000000000000200022200200200222236BCCCCCCCCBCCCCCCCCBBBAA988775543322000000000000223445678889AABBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[418] <= 3840'h5555666677777777778888888888898999A99A9A9AAAAAAAAAAAAAAAAAAABAABAAAAAAAAAABA732222220202222000200022020000020200002020000000000000022020200000000000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020002000000000000000000000200000202002000022024337BCCCCCCCCCCCCCCBCBBBA998887555332000000000000022345567888AABBBBBCBBBBBBBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB555555555555666677777777778888888888898999A99A9A9AAAAAAAAAAAAAAAAAAABAABAAAAAAAAAABA732222220202222000200022020000020200002020000000000000022020200000000000000000000000000000000000000000000000000000000000000000000000000022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020002000000000000000000000200000202002000022024337BCCCCCCCCCCCCCCBCBBBA998887555332000000000000022345567888AABBBBBCBBBBBBBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[419] <= 3840'h556666667777777778888888888998999999A9AAAAAAAAAAAAAAAAAAAAAAAAAAABABAAAABBBBA73222002022020020002020000200200000000202000000000200200222222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000022220235347BCCCCCCCCCCCCCCCBBBBA998876544322000000000000233455678899ABBBBBCBBCBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB55555555556666667777777778888888888998999999A9AAAAAAAAAAAAAAAAAAAAAAAAAAABABAAAABBBBA73222002022020020002020000200200000000202000000000200200222222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000022220235347BCCCCCCCCCCCCCCCBBBBA998876544322000000000000233455678899ABBBBBCBBCBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[420] <= 3840'h556566676777777778888888888889999999A9AAAAAAAAAAAAAAAAAAAAAAAAABAAAABABAAABBB95222202200200202002002020000002000000000200000000020202222332000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002200000000000000000200000000002002022246348CCCCCCCCCCCCCCCBBBBAA8887654432200000000000022344567888AABBBBCBBCBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB55555555556566676777777778888888888889999999A9AAAAAAAAAAAAAAAAAAAAAAAAABAAAABABAAABBB95222202200200202002002020000002000000000200000000020202222332000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002200000000000000000200000000002002022246348CCCCCCCCCCCCCCCBBBBAA8887654432200000000000022344567888AABBBBCBBCBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[421] <= 3840'h566666676777777788888888888999999999A9A9AAAAAAAAAAAAAAAAAAABAAAAABAAAAABBBBABB8422202022202000002020020020000000000000000000000002022222022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000202000000000000000000000000000200020222458558CCCCCCBCBCCCCCBBBBA99887754432200000000000022345567888AABBCBCCBBBCBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBB55555555566666676777777788888888888999999999A9A9AAAAAAAAAAAAAAAAAAABAAAAABAAAAABBBBABB8422202022202000002020020020000000000000000000000002022222022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000202000000000000000000000000000200020222458558CCCCCCBCBCCCCCBBBBA99887754432200000000000022345567888AABBCBCCBBBCBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBB;
		rom_data[422] <= 3840'h556666677777777778888888888889999999A99AAAAAAAAAAAAAAAAAAAAAAAABAAABABAAABBABBA742222220022202000020002002020000000000020000000000202022222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000022000000000000000200000000000002022023578559CCCCCCCCCCCCCBCBBAA98876554322200000000000233455678899ABBBBBBBBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBB55555555556666677777777778888888888889999999A99AAAAAAAAAAAAAAAAAAAAAAAABAAABABAAABBABBA742222220022202000020002002020000000000020000000000202022222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000022000000000000000200000000000002022023578559CCCCCCCCCCCCCBCBBAA98876554322200000000000233455678899ABBBBBBBBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBB;
		rom_data[423] <= 3840'h66566667677777777788888888889889999A99A9AAAAAAAAAAAAAAAAAAAAAAAAABAAAAABBBABABBA63220202220200020002020020200002000000000002000000002222222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000000000002000000000020202220234587469CCCCCCCCCCCCBCBBBA98877554322000000000000223455678899BBBBCCBBBBBBCBCBCBBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB5555555566566667677777777788888888889889999A99A9AAAAAAAAAAAAAAAAAAAAAAAAABAAAAABBBABABBA63220202220200020002020020200002000000000002000000002222222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000000000002000000000020202220234587469CCCCCCCCCCCCBCBBBA98877554322000000000000223455678899BBBBCCBBBBBBCBCBCBBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[424] <= 3840'h5565666667677777777878888888888999999999A9AAA9999A9AAAAAAAAAAAABAAAAABAAAABABAAB9522222020202200022020202020200002000000000000000000002020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000220000000000000200000000000000000000020000000000002022223479547BCCCCCCBCBCCCCCBBA9987764432220000000000022345567889AABBBBBBCCCCBBBBBBBCBBCBCBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB555555555565666667677777777878888888888999999999A9AAA9999A9AAAAAAAAAAAABAAAAABAAAABABAAB9522222020202200022020202020200002000000000000000000002020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000220000000000000200000000000000000000020000000000002022223479547BCCCCCCBCBCCCCCBBA9987764432220000000000022345567889AABBBBBBCCCCBBBBBBBCBBCBCBCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[425] <= 3840'h56565666767777777777888888888888999999999A999A9A9A9AAAAAAAAAAAAAABAAAAABBBBBBBBBB8522022020220002220200020220000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000002000000002000000000000000000000000000000000000000020020020222045448A9459CCCCCCCCCCCCCBBBBA988755432200000000000022344577889AABBBBCCCBBBCBBBCBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB5555556556565666767777777777888888888888999999999A999A9A9A9AAAAAAAAAAAAAABAAAAABBBBBBBBBB8522022020220002220200020220000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000002000000002000000000000000000000000000000000000000020020020222045448A9459CCCCCCCCCCCCCBBBBA988755432200000000000022344577889AABBBBCCCBBBCBBBCBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[426] <= 3840'h5555666667677777777788888888888898999999999A9A9A99A9AAAAAAAAAAABAABAABAAABBABAABBB84220022200200002002200002220000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002220028B8AEE847ACCCCCCCCCCCCCCBBA9887654422200000000000223445678899ABBBBBBBBCCBCBBCBBBBBBBCCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB555566555555666667677777777788888888888898999999999A9A9A99A9AAAAAAAAAAABAABAABAAABBABAABBB84220022200200002002200002220000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002220028B8AEE847ACCCCCCCCCCCCCCBBA9887654422200000000000223445678899ABBBBBBBBCCBCBBCBBBBBBBCCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[427] <= 3840'h55665666667777777778787888888888889899899999999A9A9AAAAA9AAAAAAAABAAAAAAAAAAABBABBB742220002202000202000202020000000002000002000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000002202027EEEEEE559CCCCCCCCCCCCCBBBAA98775442220000000000022344567889AABBBBCCBCCBBBCBBBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB5566555555665666667777777778787888888888889899899999999A9A9AAAAA9AAAAAAAABAAAAAAAAAAABBABBB742220002202000202000202020000000002000002000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000002202027EEEEEE559CCCCCCCCCCCCCBBBAA98775442220000000000022344567889AABBBBCCBCCBBBCBBBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[428] <= 3840'h55565566666677777777787888888888889898999999999999999999A9AAAAAAAAAABAABABBAAAABABAA7322222020200000000000000200000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000002000200202027EEEEEE758BCCCCBCCCCBCBCCBAA988765432200000000000023445678899ABBBCBCBCBCBCBBBBCBBBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB5665655555565566666677777777787888888888889898999999999999999999A9AAAAAAAAAABAABABBAAAABABAA7322222020200000000000000200000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000002000200202027EEEEEE758BCCCCBCCCCBCBCCBAA988765432200000000000023445678899ABBBCBCBCBCBCBBBBCBBBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[429] <= 3840'h5555565666666777777777778888888888898989998999999999A9AA99AAAAAAAABAAAAAABAAAAAAAABAA6320202000202000000200200020000000000000000000000000000000000000000000220000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000002220000000000000000000000000000000000000000000000000020203BEEEEEE758ACCCCBCCCCCCCBCBAA998765433200000000000023345678899ABBCBCCCBCBCBBBCBCBBCBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB666665565555565666666777777777778888888888898989998999999999A9AA99AAAAAAAABAAAAAABAAAAAAAABAA6320202000202000000200200020000000000000000000000000000000000000000000220000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000002220000000000000000000000000000000000000000000000000020203BEEEEEE758ACCCCBCCCCCCCBCBAA998765433200000000000023345678899ABBCBCCCBCBCBBBCBCBBCBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[430] <= 3840'h555555555566677777777777788888888988899898989889999999999999AAAAAAAAAAABAABABABABAABAA532020202000220002000002002020000000020000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002002028EEEEEA779BBCCCCCCCCCBBCCBBAA98875543220000000000023345577899ABBBCCCBBCBCBCBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB66656555555555555566677777777777788888888988899898989889999999999999AAAAAAAAAAABAABABABABAABAA532020202000220002000002002020000000020000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002002028EEEEEA779BBCCCCCCCCCBBCCBBAA98875543220000000000023345577899ABBBCCCBBCBCBCBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[431] <= 3840'h5555555565666667777777778788888888889889898989898999899999A9AAAAAAAABABAAAAABABAAAAAABA5222020202020000202000002000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000020002025CEEEC978ABCCCCCCCCCBCBCCBBBA98876543320000000000022345577899ABBBCBCBCCBCBCBBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB666555555555555565666667777777778788888888889889898989898999899999A9AAAAAAAABABAAAAABABAAAAAABA5222020202020000202000002000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000020002025CEEEC978ABCCCCCCCCCBCBCCBBBA98876543320000000000022345577899ABBBCBCBCCBCBCBBCBCBCBCBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[432] <= 3840'h55555555556566667777777778888888888898988989898888898999999A9AAAAAAAAAAABABAAAABABAAABB9622020000000200000020000220200000000000000000000000000000000000200000000000000000000000000022000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000022000000000000000000000000000000002200248ECBA99ACCCCCCCCCCCCCCCBCBBAA9877553322000000000002344577899ABBBCCCBCBCBCBCCBBBBBBBBBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB6565555555555555556566667777777778888888888898988989898888898999999A9AAAAAAAAAAABABAAAABABAAABB9622020000000200000020000220200000000000000000000000000000000000200000000000000000000000000022000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000022000000000000000000000000000000002200248ECBA99ACCCCCCCCCCCCCCCBCBBAA9877553322000000000002344577899ABBBCCCBCBCBCBCCBBBBBBBBBBBCBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[433] <= 3840'h5555555555656666667777778888888888888888888888888888988999999A9AAAAABABAAAAABAAAABABAABB95320202020200000200000000200000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000020200248CCBBBBCCCCCCCCCCCCCBCCCCBBAA9887654322000000000002344567789ABBBCCBCCCCBCBCBCBCBBCBCBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBB555555555555555555656666667777778888888888888888888888888888988999999A9AAAAABABAAAAABAAAABABAABB95320202020200000200000000200000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000020200248CCBBBBCCCCCCCCCCCCCBCCCCBBAA9887654322000000000002344567789ABBBCCBCCCCBCBCBCBCBBCBCBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBB;
		rom_data[434] <= 3840'h55555555555555656667777778888888889888888888888888888989999999AAAAAAAAAAAABAABABAAAABAABB953220200022200000000200202220000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200220248CCCCCCCCCCCCCCCCCCCCCBCBBBAA9987755332000000000002334567889ABBBCBCBBBCBCBCBCCCBCBCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBB5555555555555555555555656667777778888888889888888888888888888989999999AAAAAAAAAAAABAABABAAAABAABB953220200022200000000200202220000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200220248CCCCCCCCCCCCCCCCCCCCCBCBBBAA9987755332000000000002334567889ABBBCBCBBBCBCBCBCCCBCBCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBB;
		rom_data[435] <= 3840'h555555555555555565677777788888888888888888888888888888889999A9A9AAAAAAAAAAAAAAAAABAAAAAAAB9520202020202000000200202202200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000020000000000002000000000000000000000000000000000022222258BCCCBCCCCCCCBCBCBCBCBCCBCBAA99877654322000000000022345677899ABBCCBCBCCBCBCBCBBBBCBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB55555555555555555555555565677777788888888888888888888888888888889999A9A9AAAAAAAAAAAAAAAAABAAAAAAAB9520202020202000000200202202200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000020000000000002000000000000000000000000000000000022222258BCCCBCCCCCCCBCBCBCBCBCCBCBAA99877654322000000000022345677899ABBCCBCBCCBCBCBCBBBBCBCBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[436] <= 3840'h545555555555555556667777777888888888888888888888888888888899999AAAAAAAAAAAAABAABAAABAAAAABB9520202000002020200000022222020000200220002320000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000230000000000000000000000000000000000000000020000000022000000200000000000000000000000000000000002020025ACCCCCCBCBCCCCCCCCCCCCCCCBBBA99887655332000000000022345677889ABBBCBCBCBBCCCBCBCCCBCBCBCBCBBBCBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB55555555545555555555555556667777777888888888888888888888888888888899999AAAAAAAAAAAAABAABAAABAAAAABB9520202000002020200000022222020000200220002320000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000230000000000000000000000000000000000000000020000000022000000200000000000000000000000000000000002020025ACCCCCCBCBCCCCCCCCCCCCCCCBBBA99887655332000000000022345677889ABBBCBCBCBBCCCBCBCCCBCBCBCBCBBBCBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
		rom_data[437] <= 3840'h5454545555555555556677777787788888888888888888787888888888989999AAAAAAAAAABAAABAABAAAAABAABB85320200200020000202020222220000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000202000000000000000000000000000000000020225ACCCCCCBCBCCCCCCCCCBCBCBCBBBA99887654432000000000022344567889AABCCCBCCCBCCBBCBCBBBCBCBCBCBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBB555555445454545555555555556677777787788888888888888888787888888888989999AAAAAAAAAABAAABAABAAAAABAABB85320200200020000202020222220000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022000000202000000000000000000000000000000000020225ACCCCCCBCBCCCCCCCCCBCBCBCBBBA99887654432000000000022344567889AABCCCBCCCBCCBBCBCBBBCBCBCBCBBCBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBB;
		rom_data[438] <= 3840'h44444544455555555556677777777778788778887878777777778888888889999AAAAAAAAAAABAAAAAAAABAABABAB9630202022000220200000022222202000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022020000000000000000000000000000000000202020259CCCCCBCBCCCBCBCBCBCCCBCCCBBBA9887755432200000000022334567889AABCBCBCBCBCCBCBCBCCCCBCBCBCBCBBBCBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBB5555545444444544455555555556677777777778788778887878777777778888888889999AAAAAAAAAAABAAAAAAAABAABABAB9630202022000220200000022222202000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022020000000000000000000000000000000000202020259CCCCCBCBCCCBCBCBCBCCCBCCCBBBA9887755432200000000022334567889AABCBCBCBCBCCBCBCBCCCCBCBCBCBCBBBCBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBB;
		rom_data[439] <= 3840'h444445454545455555566667777777777777777777777777777787888889999999AAAAAAAABAAABABABABAAAAAABBB9632020200020200020000223202000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000200020236ACCCCCCCCCCBCCCCCCCCCBCCBBBBAA9987765543200000000002335567889AABBCBCCCCBCBCCCBBCBBBCBCBCCCBBCCBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABA55444444444445454545455555566667777777777777777777777777777787888889999999AAAAAAAABAAABABABABAAAAAABBB9632020200020200020000223202000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000200020236ACCCCCCCCCCBCCCCCCCCCBCCBBBBAA9987765543200000000002335567889AABBCBCCCCBCBCCCBBCBBBCBCBCCCBBCCBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABA;
		rom_data[440] <= 3840'h44344444444444555555556667777777777777777777777777777778888888899999AAAAAAAABAAAAAAAABABAAAABBAA7322220200002000020002322222020000000000000020000222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000002000202037BCCCCCCCCCBCBCBCBCBCBCCCBBBBAA98887766543200000000223345577899ABBBCBCBCBCCCBCBCCBCCCBCBCBCBCBBBCBBCCBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBB4444444444344444444444555555556667777777777777777777777777777778888888899999AAAAAAAABAAAAAAAABABAAAABBAA7322220200002000020002322222020000000000000020000222000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000002000202037BCCCCCCCCCBCBCBCBCBCBCCCBBBBAA98887766543200000000223345577899ABBBCBCBCBCCCBCBCCBCCCBCBCBCBCBBBCBBCCBCBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBB;
		rom_data[441] <= 3840'h3434334344344444555555556667677776777676666666666777777778888889999AAAAAAABAAABAAABAAAAAAAABABABB85222000200002000000023322220222000000000000020222202202000000000000000000000000000000000000000000000000000000000002000020000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000200200238CCCCCCCCCCCCCCCBCCCCCCBBBBBBAA99887777754320000000023345578899ABBCCBCCCBCBCBCBCBBCCBBCBCBCBCBCBBBCBCBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBABA544444343434334344344444555555556667677776777676666666666777777778888889999AAAAAAABAAABAAABAAAAAAAABABABB85222000200002000000023322220222000000000000020222202202000000000000000000000000000000000000000000000000000000000002000020000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000200200238CCCCCCCCCCCCCCCBCCCCCCBBBBBBAA99887777754320000000023345578899ABBCCBCCCBCBCBCBCBBCCBBCBCBCBCBCBBBCBCBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBABA;
		rom_data[442] <= 3840'h333333333343344445555555556666666666666666666566566777777888888899999AAAAAAABAAABAABABABABAAAAABBB853220200020002002002332222222220000000000002220220202202002000000000000000000000000000000000000000000000000000000000000202020000020000000000000000000000000000000000000000002002000000000000000000000000000000020000000002002002248CCCCCCCCCCCCCCBCCCCBCBCCBCBBBBAA988888875432000000022345577899ABBBCBCBCBCCCBCBCBCCBCBCBCBCBCBCBCCBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBB45443433333333333343344445555555556666666666666666666566566777777888888899999AAAAAAABAAABAABABABABAAAAABBB853220200020002002002332222222220000000000002220220202202002000000000000000000000000000000000000000000000000000000000000202020000020000000000000000000000000000000000000000002002000000000000000000000000000000020000000002002002248CCCCCCCCCCCCCCBCCCCBCBCCBCBBBBAA988888875432000000022345577899ABBBCBCBCBCCCBCBCBCCBCBCBCBCBCBCBCCBCBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBB;
		rom_data[443] <= 3840'h33333333333344445455555555555655656565655555555555566777778788889899AAAAAABABABABAAAAAABABABAAAABBB9642202020000000000023332322222220000000022020200202202002002022200002200000000000000000000000000000000200000020000200000000002000000000000000000000000000000000000000000000202000000000220000000000000000000002000000000002002238CCCCCBCCCCCCCCCCCCBCCCCBCBCBBBBAA99889987543200000002344567889ABBBCCCCCBCBCBCBCBCBBCBCBCBCBCBCBCBBCBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBABAB4444333333333333333344445455555555555655656565655555555555566777778788889899AAAAAABABABABAAAAAABABABAAAABBB9642202020000000000023332322222220000000022020200202202002002022200002200000000000000000000000000000000200000020000200000000002000000000000000000000000000000000000000000000202000000000220000000000000000000002000000000002002238CCCCCBCCCCCCCCCCCCBCCCCBCBCBBBBAA99889987543200000002344567889ABBBCCCCCBCBCBCBCBCBBCBCBCBCBCBCBCBBCBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBABAB;
		rom_data[444] <= 3840'h333233333333334444445555555555555555555555555555555666777778888888999AAAAAAAAAAAAABAABAAAAAAABAAAAABA8430202020000000022322322223222222020200222020222002220222222222222022200002200000000000000000000000000002020200000000022002000000000000000000000000000000000000020000000200000022000000000000000000000000000000000000022020248CCCCBCCCCCCCCCCCCBCCCCBCCBCCBCBBBAAA99998765200000002234567789ABBCCBCBCBCCCBCCCCCCCBBBBCBCBCBCBCBCCBCBCBBBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBABBBBB44343333333233333333334444445555555555555555555555555555555666777778888888999AAAAAAAAAAAAABAABAAAAAAABAAAAABA8430202020000000022322322223222222020200222020222002220222222222222022200002200000000000000000000000000002020200000000022002000000000000000000000000000000000000020000000200000022000000000000000000000000000000000000022020248CCCCBCCCCCCCCCCCCBCCCCBCCBCCBCBBBAAA99998765200000002234567789ABBCCBCBCBCCCBCCCCCCCBBBBCBCBCBCBCBCCBCBCBBBBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBABBBBB;
		rom_data[445] <= 3840'h3323223232333334444454555555555555555555555555555555566777778888889999AAAAAAAABAAAAABAABAABABAAABABABB95220202000002000222223333233222222220202222022222332222202222222220222220020000200000000200000000020202220020222020200020002202000000000000000000000000000000000000000200000000000000000000000000000000000000000000020002248BCCCCCCBCCCCCCBCBCCBCBCCBCCCCCCBCBBAA9AA9986430000000233557779AABBCBCCBCBCBCCCBCBCBCBCCCBCBCBCBCBCBBBBCBCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBBAAAA444333333323223232333334444454555555555555555555555555555555566777778888889999AAAAAAAABAAAAABAABAABABAAABABABB95220202000002000222223333233222222220202222022222332222202222222220222220020000200000000200000000020202220020222020200020002202000000000000000000000000000000000000000200000000000000000000000000000000000000000000020002248BCCCCCCBCCCCCCBCBCCBCBCCBCCCCCCBCBBAA9AA9986430000000233557779AABBCBCCBCBCBCCCBCBCBCBCCCBCBCBCBCBCBBBBCBCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABBBAAAA;
		rom_data[446] <= 3840'h23223222222333333444444455555555555555555555555555555567777777888898999AAAAAAAAABABAAAAABAAAAABAAABAABBA63202022020000022222223333333333332220002222022234322222222222232200322220002200000000000000000000002020220002020202222222202000000000000000000020000000000000000002000020002000000000000000000000000000000000020020220259BCBCBCBCCCBCBCBCCCCBCCCCCCCCCCCCCCBBAA9AA9875420000000234557889ABBCCCCBCBCCCCBCCCCCCCCBCBCBCBCBCBCBCBCBCBBCBBBBCBCBBBBBCBBBBBBBBBBBBBBBBBBBBBABABAAABABBAB4443332323223222222333333444444455555555555555555555555555555567777777888898999AAAAAAAAABABAAAAABAAAAABAAABAABBA63202022020000022222223333333333332220002222022234322222222222232200322220002200000000000000000000002020220002020202222222202000000000000000000020000000000000000002000020002000000000000000000000000000000000020020220259BCBCBCBCCCBCBCBCCCCBCCCCCCCCCCCCCCBBAA9AA9875420000000234557889ABBCCCCBCBCCCCBCCCCCCCCBCBCBCBCBCBCBCBCBCBBCBBBBCBCBBBBBCBBBBBBBBBBBBBBBBBBBBBABABAAABABBAB;
		rom_data[447] <= 3840'h22222222222232333334444444445555555555555555455555555566777777888889999AAAAAAABAAAAABABAAABABAAABAAAAABBA85202002020000222222222222323222222333222202223222223222223233332223222022020202000000200200000202202020202200020020220220202000000000000000002000000000202000202202000022000020200000000000000000000000000000002020036ACCBCCCCCCBCCCCCCCBCBCCBCCBCCCCCCCCCBBBA9A9976432000000223456789AABBCBBCCCCBCCCCCBCBCBCBCCBCBCCBCBCBCBCBBBCCBBCBBBBBBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABB4333323222222222222232333334444444445555555555555555455555555566777777888889999AAAAAAABAAAAABABAAABABAAABAAAAABBA85202002020000222222222222323222222333222202223222223222223233332223222022020202000000200200000202202020202200020020220220202000000000000000002000000000202000202202000022000020200000000000000000000000000000002020036ACCBCCCCCCBCCCCCCCBCBCCBCCBCCCCCCCCCBBBA9A9976432000000223456789AABBCBBCCCCBCCCCCBCBCBCBCCBCBCCBCBCBCBCBBBCCBBCBBBBBBCBCBBCBBBBBBBBBBBBBBBBBBBBBBBBABBBBBABB;
		rom_data[448] <= 3840'h322222222222232333334344444444455555555454445455555555566777777888889999AAAAAAAABABAAAAABABAAAABAABABAABBB974202020202002200000202022022022456643332222222222222232333333322322220222220202002002002202020202000000000000000202202022202020000000000000000000000002002222022020200020000000000000000000000000000000000000200236ACCCBCBCCBCCCBCBCCCCCCCCCBCCCCCCCCCBBBAAA999875320000000234557789ABBCCCCCBBCCCBCBCCCCCCCCCBCCCBCBCBCBCBCCCBCBBBBCBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABBB33333322322222222222232333334344444444455555555454445455555555566777777888889999AAAAAAAABABAAAAABABAAAABAABABAABBB974202020202002200000202022022022456643332222222222222232333333322322220222220202002002002202020202000000000000000202202022202020000000000000000000000002002222022020200020000000000000000000000000000000000000200236ACCCBCBCCBCCCBCBCCCCCCCCCBCCCCCCCCCBBBAAA999875320000000234557789ABBCCCCCBBCCCBCBCCCCCCCCCBCCCBCBCBCBCBCCCBCBBBBCBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABBB;
		rom_data[449] <= 3840'h222222222222232333333343434444445444444444444545555555556777777888889999AAAAABAAAAAABAAAAAAABABAABAAAABABBBA753202222002220020202020000020246788797322222222323333344333233323322222222222022222222220202000000000000000200000220202020220202020000202000000020202020202022020200200020000000000000000000000000000000020220237BCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCBBBBBAAA99875422000000223457788AABBCBCBCCCBCCCCCCBCBCBCBBCCCCCBCBCBCBCBBBCBBCBCBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBABABBAAAAABA33323222222222222222232333333343434444445444444444444545555555556777777888889999AAAAABAAAAAABAAAAAAABABAABAAAABABBBA753202222002220020202020000020246788797322222222323333344333233323322222222222022222222220202000000000000000200000220202020220202020000202000000020202020202022020200200020000000000000000000000000000000020220237BCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCBBBBBAAA99875422000000223457788AABBCBCBCCCBCCCCCCBCBCBCBBCCCCCBCBCBCBCBBBCBBCBCBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBABABBAAAAABA;
		rom_data[450] <= 3840'h2222222202222223233333333343443444444444444444555555555566777777888889999AAAAAAAAABAABABAABAAAAAAAAABABABABBA8532222222022220202020220202023558BEEB42323223223333334533333443322332222222220200000000000000000000000000000002020202000002220202022220020200200202022202020202020200000000000000000000000000000000000002202248BCCCBCBCBCCCCCBCBBCBCBCCCCCCBCCCCCCCBBAAA9998764320000002234567889AABBCCBCCCCCCBCCBCCCCCCCBCBCBCBCBCBCBCBCCBCCBBCBCCBBBBBCBCBCBBBBBBBBBBBBBBBBBBBAAAAAAAA9999AA333323222222222202222223233333333343443444444444444444555555555566777777888889999AAAAAAAAABAABABAABAAAAAAAAABABABABBA8532222222022220202020220202023558BEEB42323223223333334533333443322332222222220200000000000000000000000000000002020202000002220202022220020200200202022202020202020200000000000000000000000000000000000002202248BCCCBCBCBCCCCCBCBBCBCBCCCCCCBCCCCCCCBBAAA9998764320000002234567889AABBCCBCCCCCCBCCBCCCCCCCBCBCBCBCBCBCBCBCCBCCBBCBCCBBBBBCBCBCBBBBBBBBBBBBBBBBBBBAAAAAAAA9999AA;
		rom_data[451] <= 3840'h222220222222223232333333333433333333334343444555555555555666777787888999AAAAAAAAABAAAAAAABAABAABAABABAABBBABBA853322202032202020202002020024558CEEA3232233433333333334333444320222220202020200000000000000000000000000000000000202000200000020202220220002002222222022022020020200202000000000000000000000000000020002022259CCCCBCCCBCBCCCCCBCCCBCCCCCCCCCCCCCCBBBAA999987653320202223345567899ABBCBCCBCBCCCCCCCCBCBCBCCCCBCBCBCBCBCBCBCBCBBCBCBBCBBCBBBBBBBBBBBBBBBBBBBBBBBAAA999998888889933322222222220222222223232333333333433333333334343444555555555555666777787888999AAAAAAAAABAAAAAAABAABAABAABABAABBBABBA853322202032202020202002020024558CEEA3232233433333333334333444320222220202020200000000000000000000000000000000000202000200000020202220220002002222222022022020020200202000000000000000000000000000020002022259CCCCBCCCBCBCCCCCBCCCBCCCCCCCCCCCCCCBBBAA999987653320202223345567899ABBCBCCBCBCCCCCCCCBCBCBCCCCBCBCBCBCBCBCBCBCBBCBCBBCBBCBBBBBBBBBBBBBBBBBBBBBBBAAA9999988888899;
		rom_data[452] <= 3840'h22222222020222223232333333333333333333333334445555555555656677777788888999AAAAAAAAAAABABAAAAABAABAAAAABAABBABBA75432222222222202002020002035568CEE403542345543333334444544443000000000000000000000000000000000000000000020202000202200200000000200202022222202222222202022222000202000000000000000000000000000020002020225ACCCCBCBCBCCCCCCCCCBCBCBCCCCCCCCCCCBCBBAA9999876543322222334455678899BBBCBCBCCCCBCCBCBCCCCCCBCBCCCCCCBCBCBCBCBCBCBBCBCCBBBBBBCBCBBBBBBBBBBBBBBABAA99888888777777883333232222222222020222223232333333333333333333333334445555555555656677777788888999AAAAAAAAAAABABAAAAABAABAAAAABAABBABBA75432222222222202002020002035568CEE403542345543333334444544443000000000000000000000000000000000000000000020202000202200200000000200202022222202222222202022222000202000000000000000000000000000020002020225ACCCCBCBCBCCCCCCCCCBCBCBCCCCCCCCCCCBCBBAA9999876543322222334455678899BBBCBCBCCCCBCCBCBCCCCCCBCBCCCCCCBCBCBCBCBCBCBBCBCCBBBBBBCBCBBBBBBBBBBBBBBABAA9988888877777788;
		rom_data[453] <= 3840'h2222020222222222232323333333332333332333333444555555555555666777778788999A9AAAAAAABABAABABABAAAAAAAABBABAABBBBB96433222022220020202020220024578CE720355333555444433444444543000000002020202000000000000000000000000000000000002002000000000000000000202002222222222222222020002020200000020000000002000000000000020222237ACCCBCBCBCBCCCCCCCCCBCBCCCCCCCCCCCCCBBBAA9999877543322323344456677899ABBBCCCCCBBCBCCCCCCBCBCCCCCCBBCBBCBCBCCCBBCCBCCCBBBBBCBBCBBBBBBBBBBBBBAAAA99988877777666555777333232222222020222222222232323333333332333332333333444555555555555666777778788999A9AAAAAAABABAABABABAAAAAAAABBABAABBBBB96433222022220020202020220024578CE720355333555444433444444543000000002020202000000000000000000000000000000000002002000000000000000000202002222222222222222020002020200000020000000002000000000000020222237ACCCBCBCBCBCCCCCCCCCBCBCCCCCCCCCCCCCBBBAA9999877543322323344456677899ABBBCCCCCBBCBCCCCCCBCBCCCCCCBBCBBCBCBCCCBBCCBCCCBBBBBCBBCBBBBBBBBBBBBBAAAA99988877777666555777;
		rom_data[454] <= 3840'h22222220220222232223232232232232223232223333445555555555555566777777888899AAAAAABAAAAAAAAAAAAAAAABABAAAABBAABABB85322222233222020202020220225789632222453344443433223444453200002020000200000000000000000000000000000000200220002022020000000000000000002002222022220222202022020200020200000000000000000000000200220258BCCCCBCBCBCCCCCCCCCCCCBCCCCCCCCCCCBBCBBAA9999876554333333444555778889AABBBCCCBCCBCCCBCCBCCCCCBCBCBCCBCCBCBCBCBCBCBCBBCBCBBCBBBBBBBCBBBBBBBBAA989888875555555555455563333332222222220220222232223232232232232223232223333445555555555555566777777888899AAAAAABAAAAAAAAAAAAAAAABABAAAABBAABABB85322222233222020202020220225789632222453344443433223444453200002020000200000000000000000000000000000000200220002022020000000000000000002002222022220222202022020200020200000000000000000000000200220258BCCCCBCBCBCCCCCCCCCCCCBCCCCCCCCCCCBBCBBAA9999876554333333444555778889AABBBCCCBCCBCCCBCCBCCCCCBCBCBCCBCCBCBCBCBCBCBCBBCBCBBCBBBBBBBCBBBBBBBBAA98988887555555555545556;
		rom_data[455] <= 3840'h222222022022222223223223223223223232323333344555555555555555667777778888999A9AAAAAAAAAAAAAAABABBAABABBBAAABAABBBB742222202322020202202022020233323222223454333322222223443000000002020200000000000000000200000000000000000200200020200000000000000000000002002222202222022220202000020202202020000000000002020202200259BCCBCBCBCBCCCCCCCCCCCBCCCCCCCCCCCCBBBBBAAA999877554334344455566778889AABBBCCCCCCBCBCCCCCCCBCBCCCCCCBCCBCBCBCBCBCBCBCBCCBBCCBCBCBBCBBBCBBCBBA988877776554444444443455533332322222222022022222223223223223223223232323333344555555555555555667777778888999A9AAAAAAAAAAAAAAABABBAABABBBAAABAABBBB742222202322020202202022020233323222223454333322222223443000000002020200000000000000000200000000000000000200200020200000000000000000000002002222202222022220202000020202202020000000000002020202200259BCCBCBCBCBCCCCCCCCCCCBCCCCCCCCCCCCBBBBBAAA999877554334344455566778889AABBBCCCCCCBCBCCCCCCCBCBCCCCCCBCCBCBCBCBCBCBCBCBCCBBCCBCBCBBCBBBCBBCBBA9888777765544444444434555;
		rom_data[456] <= 3840'h2222222222222222222223223223222222222323334345555555555555556676777788889999AAAAAAAAABAAAABAAAAAAAABAAABBAABBAABB9533223333222020202202222202022232202222344332222222244220002000200200200000000000000000200000000000000000000000020220000000000000000000000000020220222020220202020000202000000000200000000022200037ACCCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCBBAAAA9A99887554433444556677788889AAABCBCCCCBCCCCBCCBCBCCBCCBCCCCCBCCCCCCCBCBCBCCBCBBCBBBCBCBBBBBBBBBBBAA98776555554333333333333455333333322222222222222222222223223223222222222323334345555555555555556676777788889999AAAAAAAAABAAAABAAAAAAAABAAABBAABBAABB9533223333222020202202222202022232202222344332222222244220002000200200200000000000000000200000000000000000000000020220000000000000000000000000020220222020220202020000202000000000200000000022200037ACCCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCBBAAAA9A99887554433444556677788889AAABCBCCCCBCCCCBCCBCBCCBCCBCCCCCBCCCCCCCBCBCBCCBCBBCBBBCBCBBBBBBBBBBBAA98776555554333333333333455;
		rom_data[457] <= 3840'h322222022022222223223222222222222232323333344555555555555555566777778888999AAAAAABABAAAAABABAAAABAABABABABBAAABBBB74233333432020220202202222002232222220022333222232223200020000000202000000000000002020020000000000000000200200200200200000000000000000020000202020202222220222020202000002000000000202020222200247BCCCBBCBCBCCCCCCCCCECCCCCCCCCCCCCCCBBAAAA999988876544344555677788889999AABBCCCBCCCCBCBCCBCCCCCCBCCCBCBCCCBCBCCBCBCCCBCCCBCBBCBBBBBCBCBCBBBBAA98765444443333322222223334433333232322222022022222223223222222222222232323333344555555555555555566777778888999AAAAAABABAAAAABABAAAABAABABABABBAAABBBB74233333432020220202202222002232222220022333222232223200020000000202000000000000002020020000000000000000200200200200200000000000000000020000202020202222220222020202000002000000000202020222200247BCCCBBCBCBCCCCCCCCCECCCCCCCCCCCCCCCBBAAAA999988876544344555677788889999AABBCCCBCCCCBCBCCBCCCCCCBCCCBCBCCCBCBCCBCBCCCBCCCBCBBCBBBBBCBCBCBBBBAA987654444433333222222233344;
		rom_data[458] <= 3840'h3222222022220222223223222322222222232232333445555555555555555667777788888999AAAABABAAAABAAAAABAAAABABABABABABABABB9632333343220200202002222202023222222222022223222222000220020200020020000000000020200020000002000000000002002002002200200000000000002000202000020202022202202202020202002000200202002020200202258CCCCBCCCCCCBCCBCCCCCCCCCECCECCBCCBBAAAA9999988877655444455677788899999AABBBCBBCCCBCBCBCCBCCCCBCBCCBCCCCCBCCCCCCCBCBCBCCBCBBCBCBCBCBBBBBBBCBA98875543323233332222202222333443333323222222022220222223223222322222222232232333445555555555555555667777788888999AAAABABAAAABAAAAABAAAABABABABABABABABB9632333343220200202002222202023222222222022223222222000220020200020020000000000020200020000002000000000002002002002200200000000000002000202000020202022202202202020202002000200202002020200202258CCCCBCCCCCCBCCBCCCCCCCCCECCECCBCCBBAAAA9999988877655444455677788899999AABBBCBBCCCBCBCBCCBCCCCBCBCCBCCCCCBCCCCCCCBCBCBCCBCBBCBCBCBCBBBBBBBCBA98875543323233332222202222333;
		rom_data[459] <= 3840'h3232222222022222222222222222222222223233334455555565655555555667777788888999AAAAAAAAAAAAABAAAAAAABAABABBBBBABABABBB83222333332202202022222020202222220202022022220200020200200000200020000000000002000220020000002000000000000020002002000000000000000002000002000020202022202200220220202002000200202020220202369CCCCCCCCCBCCCCBCBCCCCCCCECCECCCCBBBAA99A99988877665544455677888899AAAABABBBCBCCCBCCCCCCBCCCBCCCCCBCBCBCBCCCBCBCBCBCBCBCBBCBCBCBCBCBBCBCBCBCBA88754432222222222200000002223434333333232222222022222222222222222222222223233334455555565655555555667777788888999AAAAAAAAAAAAABAAAAAAABAABABBBBBABABABBB83222333332202202022222020202222220202022022220200020200200000200020000000000002000220020000002000000000000020002002000000000000000002000002000020202022202200220220202002000200202020220202369CCCCCCCCCBCCCCBCBCCCCCCCECCECCCCBBBAA99A99988877665544455677888899AAAABABBBCBCCCBCCCCCCBCCCBCCCCCBCBCBCBCCCBCBCBCBCBCBCBBCBCBCBCBCBBCBCBCBCBA88754432222222222200000002223;
		rom_data[460] <= 3840'h3332222222222222222232222222220222232323333455555566655555556667777778888999AAAAAABABAAAAAABBABBAABABBBABBBABABABBB952222222322200202002220222223020222202022020200020020200020200002020000000002002020020000002000000000002020002002002000000000000000002000002020002020002202202222220202020200200202022020358BCBCBBCBCCCCCCCCCCBBBBCCCCCCECCCCBBBAAA99A998877655554445567788999AAABBBBBBCCCCCBCCCCCCBCCCBCCCCCCBCBCCCCCCBCCCCCCCCCBCCBCCBCCCBCBCBCBBBBBBBBA987553322020202222000000000022444333333332222222222222222232222222220222232323333455555566655555556667777778888999AAAAAABABAAAAAABBABBAABABBBABBBABABABBB952222222322200202002220222223020222202022020200020020200020200002020000000002002020020000002000000000002020002002002000000000000000002000002020002020002202202222220202020200200202022020358BCBCBBCBCCCCCCCCCCBBBBCCCCCCECCCCBBBAAA99A998877655554445567788999AAABBBBBBCCCCCBCCCCCCBCCCBCCCCCCBCBCCCCCCBCCCCCCCCCBCCBCCBCCCBCBCBCBBBBBBBBA987553322020202222000000000022;
		rom_data[461] <= 3840'h32323222222222222232222322222222022232333344555566666655555566677777888889999AAAAAAAAABABAAAABAAABABAAABBABAABBBBBBB832000022320202202220022223422222020222020202020020202002000202200002002020202020200002000020200000000000002000200200200020000000000000000000202000002020202222220220020220002022202202247BCCBBCBCBCCCCCCCCCBBBBCCCBCCECCCCCBBAAA999999988755545444556778899AABBBBBBBBCCCCCCCCBCBCBCCBCCCCBCCCCCCBCBCBCCCCCCBBCBCCCCCBCBCBBCBCBCBCBCBBBBBA8754333220000000000000000000224434333332323222222222222232222322222222022232333344555566666655555566677777888889999AAAAAAAAABABAAAABAAABABAAABBABAABBBBBBB832000022320202202220022223422222020222020202020020202002000202200002002020202020200002000020200000000000002000200200200020000000000000000000202000002020202222220220020220002022202202247BCCBBCBCBCCCCCCCCCBBBBCCCBCCECCCCCBBAAA999999988755545444556778899AABBBBBBBBCCCCCCCCBCBCBCCBCCCCBCCCCCCBCBCBCCCCCCBBCBCCCCCBCBCBBCBCBCBCBCBBBBBA875433322000000000000000000022;
		rom_data[462] <= 3840'h33332322202222222222222222222202222232333344555666676665555666777777788889999AAAABABABABAAABBABABABABABAAABABABBABBBA4200000223222002000222224653222222222220222020200020000002020202220020202020200202020000202002000000002020020200202000000200000000000000000000002020020200220222222020202020220202002259CCCCCBCCCCCCCCCCCCCBCBBBBBBCCCECCCBBAAAA99999898765544445556788999AABBBBBBCCCCCBCBCBCCCCCCCCCCCBCCCCBCBCCCCCCCCCCCCCCBCBCBCCBCBCBBCBCBCBCBBBBBBB98653332220000000000000000000004443443333332322202222222222222222222202222232333344555666676665555666777777788889999AAAABABABABAAABBABABABABABAAABABABBABBBA4200000223222002000222224653222222222220222020200020000002020202220020202020200202020000202002000000002020020200202000000200000000000000000000002020020200220222222020202020220202002259CCCCCBCCCCCCCCCCCCCBCBBBBBBCCCECCCBBAAAA99999898765544445556788999AABBBBBBCCCCCBCBCBCCCCCCCCCCCBCCCCBCBCCCCCCCCCCCCCCBCBCBCCBCBCBBCBCBCBCBBBBBBB9865333222000000000000000000000;
		rom_data[463] <= 3840'h3333232222222222222323222222222022222333444555566777776666666777777788889999AAAAAAAABAAAABABABABAAAAAAABBAABAABABBABB7300020223320020202220249E943322222222222202000202002020202020200020202020200202200002022000200000000202000020020020200200000000000000000000002020222202022022202000200000202020202248ABCBCCCCCCCCCCCCCCCCCCCBBBBBBCCCCCCBBAAA9A9989888765544445557788999ABBBBCCCCCCCBCCCCCCCBCCBCBCCCCCCBCBCCCCCCCCCBCBCCBCBCCCCCCBCCBCCBCCBCBCBBCBCCCA9864332220000000000000000000002444443333333232222222222222323222222222022222333444555566777776666666777777788889999AAAAAAAABAAAABABABABAAAAAAABBAABAABABBABB7300020223320020202220249E943322222222222202000202002020202020200020202020200202200002022000200000000202000020020020200200000000000000000000002020222202022022202000200000202020202248ABCBCCCCCCCCCCCCCCCCCCCBBBBBBCCCCCCBBAAA9A9989888765544445557788999ABBBBCCCCCCCBCCCCCCCBCCBCBCCCCCCBCBCCCCCCCCCBCBCCBCBCCCCCCBCCBCCBCCBCBCBBCBCCCA9864332220000000000000000000002;
		rom_data[464] <= 3840'h33333323222222222222222222222022022232333445556667777776766777777778888889999AAAAABAAAABAAABAAAAABBBABAABBBABBBBBBBBB95200022022322020200027CEEE7323322222222222200020202002020202022020202020202020202020022022000200000000002020020020202000000000000000000000200020020222222222222220202020202020202469BCBCBCCCCCCCCECCECCCCCCCCBBBBBBCBCBBBAA9A9998888776555444556778889AABBBCBCBCCCCCCCCBCCBCCBCCCCBCBCCCCCCCBCCBCBBCCCCBCCCCCCCCBCCBCCBCCCBCCCBCBCBCBBB98743222200000000000000000000025444343333333323222222222222222222222022022232333445556667777776766777777778888889999AAAAABAAAABAAABAAAAABBBABAABBBABBBBBBBBB95200022022322020200027CEEE7323322222222222200020202002020202022020202020202020202020022022000200000000002020020020202000000000000000000000200020020222222222222220202020202020202469BCBCBCCCCCCCCECCECCCCCCCCBBBBBBCBCBBBAA9A9998888776555444556778889AABBBCBCBCCCCCCCCBCCBCCBCCCCBCBCCCCCCCBCCBCBBCCCCBCCCCCCCCBCCBCCBCCCBCCCBCBCBCBBB9874322220000000000000000000002;
		rom_data[465] <= 3840'h333333232222222222223222222222202222233344555567777777777777777777788888999A9AAAABAABABAABABABBBBAAABABBABBBBBBBABBABB73002202222232222248CEEEEEB5432222222220200020202202202220202020202002002020220200022202020200000000202002002002020200020000000000000000002000002002222232222220220200020200002378ACCCBCCCCCCCCECCECCCECECCCBCBBBBBBBBBAA9999998887766555444566778899ABBBCBCBCBCBCBBCBCCCBCCCCCBCCCCCCCCCCCCCCCCBCCCCCCCCBCCBCBCCCCCCBCCBCCBCBCBCBCBCBBA87532200000000000000000000000255444434333333232222222222223222222222202222233344555567777777777777777777788888999A9AAAABAABABAABABABBBBAAABABBABBBBBBBABBABB73002202222232222248CEEEEEB5432222222220200020202202202220202020202002002020220200022202020200000000202002002002020200020000000000000000002000002002222232222220220200020200002378ACCCBCCCCCCCCECCECCCECECCCBCBBBBBBBBBAA9999998887766555444566778899ABBBCBCBCBCBCBBCBCCCBCCCCCBCCCCCCCCCCCCCCCCBCCCCCCCCBCCBCBCCCCCCBCCBCCBCBCBCBCBCBBA875322000000000000000000000002;
		rom_data[466] <= 3840'h343333323222222222222232222222022022233344555667777777777777777777788888999A9AAAAAAAAAAAABABBAAAABABAAAABBABABABBABBBBA5202022002224547ACEEEEEEEC87542222220222220220220202220220202202202020202020202202002220200220000000020202002020202020000000000000000000000000000000233222222220020020020200359BCCCCCCBCCCCCCCCECCECCECCCCCCBBBBBABAAA9999998887755554544556778899AAABBBCBBBCBCCCCBCCCBCCCBCBCCBCBCBCCCCBCBCCBCCBCCCBCBCCCCCCCCCCBCBCCBCBCBCCBCBCBCBCBA98752200000000000000000000000055544434343333323222222222222232222222022022233344555667777777777777777777788888999A9AAAAAAAAAAAABABBAAAABABAAAABBABABABBABBBBA5202022002224547ACEEEEEEEC87542222220222220220220202220220202202202020202020202202002220200220000000020202002020202020000000000000000000000000000000233222222220020020020200359BCCCCCCBCCCCCCCCECCECCECCCCCCBBBBBABAAA9999998887755554544556778899AAABBBCBBBCBCCCCBCCCBCCCBCBCCBCBCBCCCCBCBCCBCCBCCCBCBCCCCCCCCCCBCBCCBCBCBCCBCBCBCBCBA987522000000000000000000000000;
		rom_data[467] <= 3840'h3433333323222222222222222222222022223333445556677777777777777777788888899999AAAAAABAAAABAABBABABAABAABABBBBBBBABBBBABBB842020222022358EEEEEEEEEEBBA9753222220202222220202202222020220222202020202020202020202020220020000202002002020202022202020200000000000000000202000023432222222020202002002257ACCCCCCCCCCCCCCCCCCCCCCECCECCCCCBBBBAA999999898887655544445556778899AAABBCCCBCCCCCBCBCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCBCBCBCBCCBCBCBCBCCBBB97530000000000000000000000000555444443433333323222222222222222222222022223333445556677777777777777777788888899999AAAAAABAAAABAABBABABAABAABABBBBBBBABBBBABBB842020222022358EEEEEEEEEEBBA9753222220202222220202202222020220222202020202020202020202020220020000202002002020202022202020200000000000000000202000023432222222020202002002257ACCCCCCCCCCCCCCCCCCCCCCECCECCCCCBBBBAA999999898887655544445556778899AAABBCCCBCCCCCBCBCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCBCBCBCBCCBCBCBCBCCBBB97530000000000000000000000000;
		rom_data[468] <= 3840'h43433333323222222322322222222022202223334455567777788888877778788888888999AAAAAAAAAABBAAAAAABABAABAABBBABABBABBABABBBBBB73020202020249EEEEEEEECAABBB98553455322222202022202202222202222222222022202020202020202002020202000020020202020202020200200000000000000000000020203532222022202020202023589BCCCCCCCCCCCCCCCCCCBCCCCCCECECCCCBBBAA99998898888765544444556678889AAABBBBCBCCCBCBCCCCCBCCBCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCBCCCCCCCCBCBCCCCBCBBCBBA85420000000000000000000000005555444443433333323222222322322222222022202223334455567777788888877778788888888999AAAAAAAAAABBAAAAAABABAABAABBBABABBABBABABBBBBB73020202020249EEEEEEEECAABBB98553455322222202022202202222202222222222022202020202020202002020202000020020202020202020200200000000000000000000020203532222022202020202023589BCCCCCCCCCCCCCCCCCCBCCCCCCECECCCCBBBAA99998898888765544444556678889AAABBBBCBCCCBCBCCCCCBCCBCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCBCCCCCCCCBCBCCCCBCBBCBBA8542000000000000000000000000;
		rom_data[469] <= 3840'h343333333323222222222232222222202022233345555677777888888788888888888899999AAAAAABABAABABBABABABBABBBBABBBBABBBBBBBBBBBBA6302022202225BEEEEEEA9BBBBBB98888BC8422223332222222222220222222020202202220202020202020202020000000022002020220222220200202000020000000000002000044200002200200200222569BBBBBBCCCCCCCCCCCCCCCBBBBBCCCCCCCBBBAAA998988888887755443445567788999ABBBCCCCCCBCCCCCCCCCCBCCCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCBCBCCCCCBCBCBCBCBCBCBA874200000000000000000000000055554444343333333323222222222232222222202022233345555677777888888788888888888899999AAAAAABABAABABBABABABBABBBBABBBBABBBBBBBBBBBBA6302022202225BEEEEEEA9BBBBBB98888BC8422223332222222222220222222020202202220202020202020202020000000022002020220222220200202000020000000000002000044200002200200200222569BBBBBBCCCCCCCCCCCCCCCBBBBBCCCCCCCBBBAAA998988888887755443445567788999ABBBCCCCCCBCCCCCCCCCCBCCCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCBCBCCCCCBCBCBCBCBCBCBA8742000000000000000000000000;
		rom_data[470] <= 3840'h44434333333323222232222222222220222223344555667777788888888888888888899999AAAAAAAAAABAAAAABAAAAAAAAABBBABABBBBABBBABBBBBB962220222022235887779BBBABBBAA98ABEC8545556655554444333332222222222222220202020202202222222220202002020200220222020202020200220000000000000000000200002002200220223568ABBAAABBBCCCCCCECCCCBCBBBBABBCCCCCBBBBA998988888877776554444566778899AABBCBCBBCBCCCCCCCBCCCBCCBCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCBCBCBCBCBCCBCBCBCBB98530000000000000000000000005555554444434333333323222232222222222220222223344555667777788888888888888888899999AAAAAAAAAABAAAAABAAAAAAAAABBBABABBBBABBBABBBBBB962220222022235887779BBBABBBAA98ABEC8545556655554444333332222222222222220202020202202222222220202002020200220222020202020200220000000000000000000200002002200220223568ABBAAABBBCCCCCCECCCCBCBBBBABBCCCCCBBBBA998988888877776554444566778899AABBCBCBBCBCCCCCCCBCCCBCCBCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCBCBCBCBCBCCBCBCBCBB9853000000000000000000000000;
		rom_data[471] <= 3840'h4444334333323223222222232222222220223334455567777888888888888888888898999AAAAAABABBAAABABAABABBABBABABABBBBABABBABBBBBBBBB973020222202223247ABBBBBBBBBAA98888878899AA9989888887775555433222222202222202202202202220200202202000220202202222220220022200220000000000000020200002002002202235799AAAAAABBBBBCCCECECCCCBBBBBAABBBBBBBAAAAA99888888887776555445556788899AABBBCCBCCBCBBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCBBA863200000000000000000000000555555444444334333323223222222232222222220223334455567777888888888888888888898999AAAAAABABBAAABABAABABBABBABABABBBBABABBABBBBBBBBB973020222202223247ABBBBBBBBBAA98888878899AA9989888887775555433222222202222202202202202220200202202000220202202222220220022200220000000000000020200002002002202235799AAAAAABBBBBCCCECECCCCBBBBBAABBBBBBBAAAAA99888888887776555445556788899AABBBCCBCCBCBBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCBBA863200000000000000000000000;
		rom_data[472] <= 3840'h4444433333332322322232222222220222222334455567778888888888888888889899999AAAAAAABAABBBAAAABAAAABAABABBBBBABBBBBBBABABBBBBBBA743202022223358ABBBBBBBBABBBAA999999AABABBBABABAAAA9988888765555544322222202202002202022222002020202022202222222333222220220200000000000000000000002002022345689AA999AA9AABBBBCCCECCCCCCCBBBBBAAAAAAA99999898888888776655545556777889AAABBBBBBCCBCCCBCCCCCBBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBBCCBCBCBCCBCBB874300000000000000000000000555555554444433333332322322232222222220222222334455567778888888888888888889899999AAAAAAABAABBBAAAABAAAABAABABBBBBABBBBBBBABABBBBBBBA743202022223358ABBBBBBBBABBBAA999999AABABBBABABAAAA9988888765555544322222202202002202022222002020202022202222222333222220220200000000000000000000002002022345689AA999AA9AABBBBCCCECCCCCCCBBBBBAAAAAAA99999898888888776655545556777889AAABBBBBBCCBCCCBCCCCCBBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBBCCBCBCBCCBCBB874300000000000000000000000;
		rom_data[473] <= 3840'h44443434333332232222222232222222222233345556677888888898988988888998999AAAAAAAAAABAAAABBBBABABBABAAABBBABBBABBABABBBBBBBBBBBA8754333344579BBBBBBBBBBBABBBBBAAABABBBABBBBBBBBBAABAABBAA9999988887765444432222220202202020202222222333432233349BBA853322220200200000000202020000002223457788999999A99A99AABBBCCCCECCCCCCCBBAAA9A9989989888888888776555545556778889AAABBBCBCCBCCBBCBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCCBCBCBCCCB9875333202000000000000000006555555544443434333332232222222232222222222233345556677888888898988988888998999AAAAAAAAAABAAAABBBBABABBABAAABBBABBBABBABABBBBBBBBBBBA8754333344579BBBBBBBBBBBABBBBBAAABABBBABBBBBBBBBAABAABBAA9999988887765444432222220202202020202222222333432233349BBA853322220200200000000202020000002223457788999999A99A99AABBBCCCCECCCCCCCBBAAA9A9989989888888888776555545556778889AAABBBCBCCBCCBBCBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCCBCBCBCCCB987533320200000000000000000;
		rom_data[474] <= 3840'h544444343333323232322232222222222222334445567778888889999989899998999999AAAAABABAABABAAAAAAABAABBBBABABBBABBABBBBBBBBBBBBBBBBBA98767789AACBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBABBBAABABBBABABBABBABAA9988877655544333333322333344334567775433236EEEEEC7543222222220220202000020222234567789999999999A9A9999BBBBBCCCCCCECCCCCBBAAA9988898888888887775554545557778899AABBBCBCBCBCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCCCBCBBA9876555544444330000000002266655555544444343333323232322232222222222222334445567778888889999989899998999999AAAAABABAABABAAAAAAABAABBBBABABBBABBABBBBBBBBBBBBBBBBBA98767789AACBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBABBBAABABBBABABBABBABAA9988877655544333333322333344334567775433236EEEEEC7543222222220220202000020222234567789999999999A9A9999BBBBBCCCCCCECCCCCBBAAA9988898888888887775554545557778899AABBBCBCBCBCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCCCBCBBA98765555444443300000000022;
		rom_data[475] <= 3840'h55444343333333232222222232322222222333345556777888999999999999989999A9AAAAABAAAAAAAAABABAAAABBBBABABBBABBBBBBBABABABBABABABBBBBBBBAAABBBBBBBBBABBBBBBBBABBBABABABBBBABABAABBAABBBBBABABBBBBBBBBBBBBBBBAAA998887667776557777888889AABB9854224BEEEEE94543343343222020222333334455667888899898899999999999AAAABBBCCCCCCCCBBBBAA999889998888777776555444556778889AAABBCCBCBCBCBCCCCCCBCCCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCCBBAA9888777677553320000022326666555555444343333333232222222232322222222333345556777888999999999999989999A9AAAAABAAAAAAAAABABAAAABBBBABABBBABBBBBBBABABABBABABABBBBBBBBAAABBBBBBBBBABBBBBBBBABBBABABABBBBABABAABBAABBBBBABABBBBBBBBBBBBBBBBAAA998887667776557777888889AABB9854224BEEEEE94543343343222020222333334455667888899898899999999999AAAABBBCCCCCCCCBBBBAA999889998888777776555444556778889AAABBCCBCBCBCBCCCCCCBCCCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCCBBAA988877767755332000002232;
		rom_data[476] <= 3840'h554444434333333333232232322232222223334455567778898999999999999999A9AAAAAAAAABABABABAABABABABABBBBABABBBABABABABBBBBBBABABBBBBBBBCBBBCBBBBBBBBBABBBABBBBBABBABBABBBBABBABBBABBBBBABBBBBBBBBBBBBBBBBBBBCBCCCBBBAAAABAA99ABBBBBBBBCCBCCCB974325AEEEE63443334554222223345667777778888888889898989999898889999AAABBBBBBBBBABABBAAA999999888877765554454556778899AABBBBBBCCBCBBCCBBCBCCCCCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCBCBBBBAAA9999887543222022233366666555554444434333333333232232322232222223334455567778898999999999999999A9AAAAAAAAABABABABAABABABABABBBBABABBBABABABABBBBBBBABABBBBBBBBCBBBCBBBBBBBBBABBBABBBBBABBABBABBBBABBABBBABBBBBABBBBBBBBBBBBBBBBBBBBCBCCCBBBAAAABAA99ABBBBBBBBCCBCCCB974325AEEEE63443334554222223345667777778888888889898989999898889999AAABBBBBBBBBABABBAAA999999888877765554454556778899AABBBBBBCCBCBBCCBBCBCCCCCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCBCBBBBAAA99998875432220222333;
		rom_data[477] <= 3840'h555444444343333323223222323222222333334555577788899999999999A99999AAAAAAAAAAAAAAAABAABAABBBABBBABAAABBABBBBBBBBBBBABBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBABBBABABBABABBBBBBBBABABBABBABBBBBBBBBBBBBBBBBBABCBCBBCBCBBBCCCBCBBCBCBBBCBCCCA854236BC833432223333222234589A9999988888888898989899898898888888899AAAAAAABBAAAAAAAAA99999988877655554444556778899AABBCBCBCCBCBCCBCCCCCCCCCCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCBCBCCCBBBBCBBBAA987553322233333366666665555444444343333323223222323222222333334555577788899999999999A99999AAAAAAAAAAAAAAAABAABAABBBABBBABAAABBABBBBBBBBBBBABBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBABBBABABBABABBBBBBBBABABBABBABBBBBBBBBBBBBBBBBBABCBCBBCBCBBBCCCBCBBCBCBBBCBCCCA854236BC833432223333222234589A9999988888888898989899898898888888899AAAAAAABBAAAAAAAAA99999988877655554444556778899AABBCBCBCCBCBCCBCCCCCCCCCCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCBCBCCCBBBBCBBBAA9875533222333333;
		rom_data[478] <= 3840'h55555444443433333323223232233232323334455567788889999A9A9A9A9AA9AAAAAAAABABABABABAAAAABBAABBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBBABBBABBABBBABBBBABABABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCBBBBCB975334432322222022222345789998888888888888989998989888888888989889AA9A9999AA9999AAAA9999988877555444444557788899AABBCBCCCBCCBCBBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCBCBCBCCCBBAA87654433233334336666665655555444443433333323223232233232323334455567788889999A9A9A9A9AA9AAAAAAAABABABABABAAAAABBAABBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBBABBBABBABBBABBBBABABABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCBBBBCB975334432322222022222345789998888888888888989998989888888888989889AA9A9999AA9999AAAA9999988877555444444557788899AABBCBCCCBCCBCBBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCBCBCBCCCBBAA8765443323333433;
		rom_data[479] <= 3840'h55555444434433333232322232322323233334555567788899999A9A9A9A9A9AAAAAAAABAAABAAAAABABABBAABAABBBABAAABBABABABABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBABBABBBABBBBBBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCBBBCBBBCBB9864332222222222334568888888888888899999999998989888888888888888989988888889999AA9999888877655444445557788899ABBBCCCBCBCBCCBCCBCBCCCBCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCBCCBBAA9876544333333443436676666655555444434433333232322232322323233334555567788899999A9A9A9A9A9AAAAAAAABAAABAAAAABABABBAABAABBBABAAABBABABABABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBBBBBABBABBBABBBBBBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCBBBCBBBCBB9864332222222222334568888888888888899999999998989888888888888888989988888889999AA9999888877655444445557788899ABBBCCCBCBCBCCBCCBCBCCCBCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCBCCBBAA987654433333344343;
		rom_data[480] <= 3840'h655555444444443333232323232323232333445555777888899A9A9A9A9AAAAAAAAAAAAAABAAAABAABABAABBAABABABBBAAABBBBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBABBBABBBBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBCBCCBBBA87655433334556778889888888888999999999999999888888888998888888888777888888899999988887765544434556678899AABBBBCCCCBCCCBCCBCCBCBBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCBBBA9887554333334444433366767666655555444444443333232323232323232333445555777888899A9A9A9A9AAAAAAAAAAAAAABAAAABAABABAABBAABABABBBAAABBBBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABBABBBABBBBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBCBCCBBBA87655433334556778889888888888999999999999999888888888998888888888777888888899999988887765544434556678899AABBBBCCCCBCCCBCCBCCBCBBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCBBBA98875543333344444333;
		rom_data[481] <= 3840'h6555554544444333333232232323232323344455567788889999AAAAAAAAAAAAAAAAAAAAAABABAABAABAABBABABABBBAAABABABABBBBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBABBBABABBBBBBBBABBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCBBBCBBBBBBBBBCBBCBBA9877778889AA9988888788888999999999999999988888888999888878888777777887788999988777755544444555778899AABBBCCBBCBCBCBCBCCBCCCCCCCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCBBBA9887755433334444433333677676766555554544444333333232232323232323344455567788889999AAAAAAAAAAAAAAAAAAAAAABABAABAABAABBABABABBBAAABABABABBBBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBABBBABABBBBBBBBABBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCBBBCBBBBBBBBBCBBCBBA9877778889AA9988888788888999999999999999988888888999888878888777777887788999988777755544444555778899AABBBCCBBCBCBCBCBCCBCCCCCCCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCBBBA9887755433334444433333;
		rom_data[482] <= 3840'h665555544444444333332332323232333334455566778888999999A9AAAAAAAAAAAAAABABAAAABAAABAABABAABABBBABBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBABBBBBABBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBCBCBCBCBCBBBCBBBBBBABBBBBBAA988888888888999999999A9999998888888899888877777666666777777788998877765544444556778899AABBBCBCCCBCCCBCCCCBCCBCBCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBA99887655433434444343332276767777665555544444444333332332323232333334455566778888999999A9AAAAAAAAAAAAAABABAAAABAAABAABABAABABBBABBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBABBBBBABBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBCBCBCBCBCBBBCBBBBBBABBBBBBAA988888888888999999999A9999998888888899888877777666666777777788998877765544444556778899AABBBCBCCCBCCCBCCCCBCCBCBCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBA998876554334344443433322;
		rom_data[483] <= 3840'h665555554444444343333232323323333344555567778889999A9A9AAAAAAAAAABAAABABABAAAAABAABBABABBBBBABBBBABAABBBBBBBABBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBABABBBBBBBBBBBBABABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBBBBBBBCBCBBBCCCCBCCCCCBBAAA98888888889999A9A999999999988888888888877555555555555666777888888776554444556678899AAABBBCCCBCBCCBCBCBBCCBCBCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBA9987765554444444443333322266667676665555554444444343333232323323333344555567778889999A9A9AAAAAAAAAABAAABABABAAAAABAABBABABBBBBABBBBABAABBBBBBBABBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBABABBBBBBBBBBBBABABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBBBBBBBCBCBBBCCCCBCCCCCBBAAA98888888889999A9A999999999988888888888877555555555555666777888888776554444556678899AAABBBCCCBCBCCBCBCBBCCBCBCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBA99877655544444444433333222;
		rom_data[484] <= 3840'h7665555554444443433333332332333334445556777888889999A9AAAAAAAAAAAAAAAAAAAAABABAAABAABAAAAABABBBABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBABBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBBCBBBCBCBCBCBCBCBBBAA9999998888899999899899999988887887777776555555454555555556778888877655545556677889AAABBBCBCBCCCBCBCBCBCBCBCBCBCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAA9988775554444445444333322220676676777665555554444443433333332332333334445556777888889999A9AAAAAAAAAAAAAAAAAAAAABABAAABAABAAAAABABBBABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBABBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBBCBBBCBCBCBCBCBCBBBAA9999998888899999899899999988887887777776555555454555555556778888877655545556677889AAABBBCBCBCCCBCBCBCBCBCBCBCBCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAA9988775554444445444333322220;
		rom_data[485] <= 3840'h7666555555444444433333233323333344455556777888899999A9AAAAAAAAAAAAABABAAAAAAAAABABABABBBBBBBAABBBABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBABABABBBBBBBBBBBBBABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBBBBCBCBCBCBCBBBCBCBCBCBCBBBBAAAAA99999999999988888889888777777776765555554454444444445567788877665555556778899ABBBBCCBCBCBCBCBCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAAA998877655454455555444333222000676777767666555555444444433333233323333344455556777888899999A9AAAAAAAAAAAAABABAAAAAAAAABABABABBBBBBBAABBBABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBABABABBBBBBBBBBBBBABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBBBBCBCBCBCBCBBBCBCBCBCBCBBBBAAAAA99999999999988888889888777777776765555554454444444445567788877665555556778899ABBBBCCBCBCBCBCBCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAAA998877655454455555444333222000;
		rom_data[486] <= 3840'h777665555545444434433333233333334455566777888889999A9A9AAAAAAAABAAAAAABABABABABABABBBBABABBBBBAABBBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBCBCBCBCBCBBCBCBCBCCBBBCBCBBCBBBBBBBBBAAAAA9A9AA9999898888888777777776665555555555554444343445578887766655567788899AABBBCCCCCCCCCCCCBCBCBCBBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBA99988777654544444455554332222020066776777777665555545444434433333233333334455566777888889999A9A9AAAAAAAABAAAAAABABABABABABABBBBABABBBBBAABBBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBCBCBCBCBCBBCBCBCBCCBBBCBCBBCBBBBBBBBBAAAAA9A9AA9999898888888777777776665555555555554444343445578887766655567788899AABBBCCCCCCCCCCCCBCBCBCBBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBA999887776545444444555543322220200;
		rom_data[487] <= 3840'h7776655555454444443433333333334445555667778888899999A9AAAAAAAABAAAABABAAAABAABAABBBABABBBBABAABBABABAABBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBABABBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCCBCBBBBBCBCCBCBCBCBBBBCBCBCBBCCCBCBBBBBBBAAAAAAAAAA999999998888777777766555566665555444333333446777766665667788999AABBBCCCCBBCBCBCCCCCBCBCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCECCCCCCCCECCECCECCCCCCCCCCCCBBAAA99988777555544443444555543332202000676677777776655555454444443433333333334445555667778888899999A9AAAAAAAABAAAABABAAAABAABAABBBABABBBBABAABBABABAABBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBABBBBABABBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCCBCBBBBBCBCCBCBCBCBBBBCBCBCBBCCCBCBBBBBBBAAAAAAAAAA999999998888777777766555566665555444333333446777766665667788999AABBBCCCCBBCBCBCCCCCBCBCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCECCCCCCCCECCECCECCCCCCCCCCCCBBAAA99988777555544443444555543332202000;
		rom_data[488] <= 3840'h7777665555544444443433333333434445556677778888889999A9AAAAAAAAAAAAABAAAAAAABAAABAABABBBABABBBBABBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCBCCCCCBCBCBCBCBCBCBCCBCBBCBBCBCCBCBBBBBBBBBAAABAABAAA9AA999887877777777666777665555433322233456777666667788899AABBBBCBCCCCCCCCCCBCBCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBA99888877655545444333344555443322020000667767777777665555544444443433333333434445556677778888889999A9AAAAAAAAAAAAABAAAAAAABAAABAABABBBABABBBBABBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCBCCCCCBCBCBCBCBCBCBCCBCBBCBBCBCCBCBBBBBBBBBAAABAABAAA9AA999887877777777666777665555433322233456777666667788899AABBBBCBCCCCCCCCCCBCBCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBA99888877655545444333344555443322020000;
		rom_data[489] <= 3840'h776666655555444444443433333344455556677778888899999A9A9AAAAAAAAAAAAABABAAABABBBABBBBBABBBBBABABABABABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBABBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCCBCBCBBBBBCBBCBCBCBCBCBCBCBCBCBCBBBBCBCCCBCBBBBBBBBBBBBBBAABA9998888787877777776665554443322222334566666677888899AABBBCCBCCCCCBCBCCCCCCCCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECECECCCCCCCCCCCCCCCCCBBAAA98887776555544444333333445554322200000066767777776666655555444444443433333344455556677778888899999A9A9AAAAAAAAAAAAABABAAABABBBABBBBBABBBBBABABABABABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBABBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCCBCBCBBBBBCBBCBCBCBCBCBCBCBCBCBCBBBBCBCCCBCBBBBBBBBBBBBBBAABA9998888787877777776665554443322222334566666677888899AABBBCCBCCCCCBCBCCCCCCCCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECECECCCCCCCCCCCCCCCCCBBAAA988877765555444443333334455543222000000;
		rom_data[490] <= 3840'h7777666555554544444434333334444555566777788888999999A9AAAAAAAAAABAAAAAAABAAAAAAABABABBBABABABBBBAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBABBBBABABBBBBBBBBBBBBBBBBABABBBBBBBBBBBBBBBBBBBBCBCBBBBBBCBCBCBCCCBCBCBCBCBCBCBCBCBCBCBCBBCBCBCBBCCCCBCBBCBBBBBBBBBBBBAA99988888877776655555443332220223345555567788889AAABBBCBCCCBCBCCCCCCBCCBCBCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCCCCCCCCCCCCECCECCECCCCCCBBBBA998877665555544443333222234455443220200023676776777777666555554544444434333334444555566777788888999999A9AAAAAAAAAABAAAAAAABAAAAAAABABABBBABABABBBBAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBABBBBABABBBBBBBBBBBBBBBBBABABBBBBBBBBBBBBBBBBBBBCBCBBBBBBCBCBCBCCCBCBCBCBCBCBCBCBCBCBCBCBBCBCBCBBCCCCBCBBCBBBBBBBBBBBBAA99988888877776655555443332220223345555567788889AAABBBCBCCCBCBCCCCCCBCCBCBCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCCCCCCCCCCCCECCECCECCCCCCBBBBA998877665555544443333222234455443220200023;
		rom_data[491] <= 3840'h77776765555554444444443443444555555677777888899999A9A9AAAAAAAAAAAABAABABABBBABABABBBBABBBABBBABBBBBABBBABABBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCCBBBCBBCBBCBCBCBCBCBCBCBCBCBCBCBBCBBCBCBCCBBCBCBCBCCBCBCBCBCBBBAAA99888877756555554433322202222334555556778899AABBBCCCCCCCCCCCBCCBCCCCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECECCCCCCCCCCCCBBBAA998876665555444433332222022233444332200223456677777777776765555554444444443443444555555677777888899999A9A9AAAAAAAAAAAABAABABABBBABABABBBBABBBABBBABBBBBABBBABABBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCCBBBCBBCBBCBCBCBCBCBCBCBCBCBCBCBBCBBCBCBCCBBCBCBCBCCBCBCBCBCBBBAAA99888877756555554433322202222334555556778899AABBBCCCCCCCCCCCBCCBCCCCCCCBCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECECCCCCCCCCCCCBBBAA99887666555544443333222202223344433220022345;
		rom_data[492] <= 3840'h777777665555544444444444444445555666777888888899999A9AAAAAAAAAAAAAAAAAAAAAAABABABBBABBBABBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCCCCBCBCBCBCCBCBCBBBCCCCCCCBCBBBBA99988877665555544433222222222335455555577899ABBBBCBCBCCCCBCBCCCCCCCCBCCBCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECCECCECCECCCCCCCCCCCCCCCBBAA9988877655555444333322222000002233343220223456767677677777777665555544444444444444445555666777888888899999A9AAAAAAAAAAAAAAAAAAAAAAABABABBBABBBABBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCCCCBCBCBCBCCBCBCBBBCCCCCCCBCBBBBA99988877665555544433222222222335455555577899ABBBBCBCBCCCCBCBCCCCCCCCBCCBCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECCECCECCECCCCCCCCCCCCCCCBBAA99888776555554443333222220000022333432202234567;
		rom_data[493] <= 3840'h77777766655545454545544444445555666777888888899999A9AAAAAAAAAAAAAAAABABAAABAAABBABABBABBBABBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBBCBCBCBCBCBCBCBCBCBCBCBCBCCBBBBBA9988887765555454333222202223344555555556789AABBCCCBCCCCCBCCCCBCBCCBCCCBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECECECCCCCBBAAA98887776555544433332222200000000022333332234567897767677777777766655545454545544444445555666777888888899999A9AAAAAAAAAAAAAAAABABAAABAAABBABABBABBBABBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBBCBCBCBCBCBCBCBCBCBCBCBCBCCBBBBBA9988887765555454333222202223344555555556789AABBCCCBCCCCCBCCCCBCBCCBCCCBCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECECECCCCCBBAAA9888777655554443333222220000000002233333223456789;
		rom_data[494] <= 3840'h777777766555554544555544445455556677777888889899999A99AAAAAAAAAAAAABABAAAAAABBABBBBBBBBABABBBBBBBBBBBBABBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCCBCCCBCBCCCBCCCCCCCCCCCCCCCCBBBAA9988877655544433332220222233445555555555789ABBBCBCCCBCBCCCCBCCCCBCCCBCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECCCECCCCCCCCCCCCCBBAA99888776555554433332222220000000000000233234456789AB67676777777777766555554544555544445455556677777888889899999A99AAAAAAAAAAAAABABAAAAAABBABBBBBBBBABABBBBBBBBBBBBABBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCCBCCCBCBCCCBCCCCCCCCCCCCCCCCBBBAA9988877655544433332220222233445555555555789ABBBCBCCCBCBCCCCBCCCCBCCCBCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECCCECCCCCCCCCCCCCBBAA99888776555554433332222220000000000000233234456789AB;
		rom_data[495] <= 3840'h7777777666555554545555555555555567777888888989999A99A9AAAAAAAAAAAAAAAAABAABBABBBABABABBBAABABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCCBBCBCBCBCCCCCBCBCBCBCBCBBBBCBCBCCBCBCBCBCBCBCBBCBBCBBCCCBCBBBBAA9988776655444333222222222334455677655455679ABCCCCCBCCCCCCCCCCBCCCCBCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCCECECCCCCCCBAAA98887776555544433332222020000000000000002223456789ABBB767677777777777666555554545555555555555567777888888989999A99A9AAAAAAAAAAAAAAAAABAABBABBBABABABBBAABABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCCBBCBCBCBCCCCCBCBCBCBCBCBBBBCBCBCCBCBCBCBCBCBCBBCBBCBBCCCBCBBBBAA9988776655444333222222222334455677655455679ABCCCCCBCCCCCCCCCCBCCCCBCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCCECECCCCCCCBAAA98887776555544433332222020000000000000002223456789ABBB;
		rom_data[496] <= 3840'h777777776655554555555555545555566777888888889999999A9A9AAAAAAAAAAABAAAAAABAAABABABBBBBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBCCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCCCBCCBCCBCCCBCCBBBBAA998887765544433332202022333455667777755455789BCCCBCCCCCCCCCCCCCCCBCCCBCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCCCCCCCBAAA998877765555544433322222200000000000000000000245789ABBCCC67777777777777776655554555555555545555566777888888889999999A9A9AAAAAAAAAAABAAAAAABAAABABABBBBBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBCCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCCCBCCBCCBCCCBCCBBBBAA998887765544433332202022333455667777755455789BCCCBCCCCCCCCCCCCCCCBCCCBCCCBCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCCCCCCCBAAA998877765555544433322222200000000000000000000245789ABBCCC;
		rom_data[497] <= 3840'h77777777665555555555555555555566777778888889999999A9A9A9AAAAAAAAAAAABABAAABBBABBBAABBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBCBCBCBCCBCBCBCBCCCCCCCCCBCBCCBCBCCCCCCCBCBCCCBCCBCCBCCCBCBBAAA998877665544333222202223334555778888775545689BBCCCCCCCCCCCCCCCCCCCCCCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCECCCCCCCCCBBBAA99988877655555443333222200000000000000000000000035789ABCCCCC7667677777777777665555555555555555555566777778888889999999A9A9A9AAAAAAAAAAAABABAAABBBABBBAABBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBCBCBCBCCBCBCBCBCCCCCCCCCBCBCCBCBCCCCCCCBCBCCCBCCBCCBCCCBCBBAAA998877665544333222202223334555778888775545689BBCCCCCCCCCCCCCCCCCCCCCCCCBCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCECCCCCCCCCBBBAA99988877655555443333222200000000000000000000000035789ABCCCCC;
		rom_data[498] <= 3840'h777777776655555555555555555556667778888888898999999A9A9A9AAAAAAAAAABABAABAAABBBABABABABBABBABBBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBCBCBCBCBCBCBCBCCCBCBCBCBBBCBBCBCCBBCCBCCBCBBCBCBCBBCCCCCCCCCCCBCBBAA9988877555443332220222233445567788899875544579BBCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECCCCCECCCCCCBBAA9998887776555554433332222000000000000000000000000024689BCCCCCCC67677677777777776655555555555555555556667778888888898999999A9A9A9AAAAAAAAAABABAABAAABBBABABABABBABBABBBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBCBCBCBCBCBCBCBCCCBCBCBCBBBCBBCBCCBBCCBCCBCBBCBCBCBBCCCCCCCCCCCBCBBAA9988877555443332220222233445567788899875544579BBCCCCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCECCCCCECCCCCCBBAA9998887776555554433332222000000000000000000000000024689BCCCCCCC;
		rom_data[499] <= 3840'h777777776655555555555555555556677778888888989999999A9A9A9AAAAAAAAAAAAAABABABBBBBABABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBCBBBCBBBCBBBCBCBCBCBCBCBCCCCBCBCBCCCCCBCCBCBCBCCBCBCCBCCCCBCCCCBCBCCBCCBBBCBBAAA98887665544332222022223344556778899A9987544578ABCBCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECECCCCCBBAA998887777655554444333222200000000000000000023333200023579ACCCCCCCC67677777777777776655555555555555555556677778888888989999999A9A9A9AAAAAAAAAAAAAABABABBBBBABABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBCBBBCBBBCBBBCBCBCBCBCBCBCCCCBCBCBCCCCCBCCBCBCBCCBCBCCBCCCCBCCCCBCBCCBCCBBBCBBAAA98887665544332222022223344556778899A9987544578ABCBCCCCCCCCCCCCCCCCCCCCCCCCCCBCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECECCCCCBBAA998887777655554444333222200000000000000000023333200023579ACCCCCCCC;
		rom_data[500] <= 3840'h7777777776655555555556666565667777888888888999999999A9A9AAAAAAAAAABAABAAAAAAABABBABBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBCCCBCBCCCCCCCBBCBCCBCCCBCBCCCCCBCCCBCCBCBCCCCBCCBCCCCBBBAA98887765554333220222233345557788899AABA975445589BBCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCCBBA99888776655555444433332222000000000000000223445666654444678ACCCCCCCCC666777777777777776655555555556666565667777888888888999999999A9A9AAAAAAAAAABAABAAAAAAABABBABBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBCCCBCBCCCCCCCBBCBCCBCCCBCBCCCCCBCCCBCCBCBCCCCBCCBCCCCBBBAA98887765554333220222233345557788899AABA975445589BBCCCCCCCCCCCCCCCCCCCCCCCBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCCBBA99888776655555444433332222000000000000000223445666654444678ACCCCCCCCC;
		rom_data[501] <= 3840'h777777777765555555566666666666777888888889999899999999A9AAAAAAAAAAAABAABAABBBBBABBBABBABABBBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBBCBCBCBCBCCBCCBCBBCBCCCCBCCBCBCCCBCBBCCCCCCCBCCCCBCCCCCCCBCBBBAA9988776554433222020222335556778899AABBBBA87544579BBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCCECCCCCCBAA988877665555544433332222020000000000000022455667889888877789ABCCCCCCCCC67777777777777777765555555566666666666777888888889999899999999A9AAAAAAAAAAAABAABAABBBBBABBBABBABABBBBABBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBBCBCBCBCBCCBCCBCBBCBCCCCBCCBCBCCCBCBBCCCCCCCBCCCCBCCCCCCCBCBBBAA9988776554433222020222335556778899AABBBBA87544579BBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCECCCECCCCCCBAA988877665555544433332222020000000000000022455667889888877789ABCCCCCCCCC;
		rom_data[502] <= 3840'h7777777777665555556667676666777778888888989899999999A99A9AAAAAAAAABAAAAAABABBBBBBBABABBBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBBBCBBBBBCBCBCBCBCBCBCBCCCCCBCCBCBCCBCCCBCBCBCCCBCBCBCCCCBCCCCCBCBCCBBAAA9988777554333220202222344556678899AAABBCCB98544568ABBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBAAA9888776655554443333222202000000000000002235567899AAABBBBA9A9ABBCCCCCCCCCC666677777777777777665555556667676666777778888888989899999999A99A9AAAAAAAAABAAAAAABABBBBBBBABABBBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBBBCBBBBBCBCBCBCBCBCBCBCCCCCBCCBCBCCBCCCBCBCBCCCBCBCBCCCCBCCCCCBCBCCBBAAA9988777554333220202222344556678899AAABBCCB98544568ABBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBAAA9888776655554443333222202000000000000002235567899AAABBBBA9A9ABBCCCCCCCCCC;
		rom_data[503] <= 3840'h777777777766555556666677776667778888889889989999999999A9AAAAAAAAAAAABABAAAABBBAABBBBBBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBCBCBCBCCBCCBCBCBCCBCCBCBCCBCBCCCCCBCBCCCCCCBCBCCBCBCCCCCBCBAA998877655443322202022334455677889AAABBBCCCCA97544589BBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBAAA9988877755554443332222202000000000000000234577899ABBBCCCCCCCCBCCCCCCCCCCCCCC76777777777777777766555556666677776667778888889889989999999999A9AAAAAAAAAAAABABAAAABBBAABBBBBBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBCBCBCBCCBCCBCBCBCCBCCBCBCCBCBCCCCCBCBCCCCCCBCBCCBCBCCCCCBCBAA998877655443322202022334455677889AAABBBCCCCA97544589BBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBAAA9988877755554443332222202000000000000000234577899ABBBCCCCCCCCBCCCCCCCCCCCCCC;
		rom_data[504] <= 3840'h777777777766655555677777777777778888888899898999999A9A9A9AAAAAAAAABAAAAABABBABBBBABBABBABBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBCBCBBBCBCCCCCCBCCCCCCBCCBCCCCBCCCBCBBCBCBCCCCBCCCCCCCCCBCCBCBBAA998887655443322020222334455677899AAABBCCCCCCBA8644579BBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAA998887777555544433322222000000000000000234556788AABCCCCCCCCCCCCCCCCCCCCCCCCCCCC67777777777777777766655555677777777777778888888899898999999A9A9A9AAAAAAAAABAAAAABABBABBBBABBABBABBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBCBCBBBCBCCCCCCBCCCCCCBCCBCCCCBCCCBCBBCBCBCCCCBCCCCCCCCCBCCBCBBAA998887655443322020222334455677899AAABBCCCCCCBA8644579BBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAA998887777555544433322222000000000000000234556788AABCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
		rom_data[505] <= 3840'h77777777777666565667777777777777888888989898999999999A9A9AAAAAAAAAAABAAAAABBBBABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBBBCCCCCBCBCBCBCBCBCCCBCCBCBCCBCCCCCBCCCCBCCCCBCCBCBCBCCBCBBBAA99887665443322020222334455777889AABBCBCCCCCCCB97545789BCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCBBAA988877777555544433322220200000000000002345567899ABBBCCCCCCCCCCCCCCCCCCCCCCCCCCCCC7767777777777777777666565667777777777777888888989898999999999A9A9AAAAAAAAAAABAAAAABBBBABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBBBCCCCCBCBCBCBCBCBCCCBCCBCBCCBCCCCCBCCCCBCCCCBCCBCBCBCCBCBBBAA99887665443322020222334455777889AABBCBCCCCCCCB97545789BCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCECCCCCCBBAA988877777555544433322220200000000000002345567899ABBBCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
		rom_data[506] <= 3840'h777777777776656666777777777777788888888898989899999999A9A9A9AAAAAABAABABAAABABBABABBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBBBCBCCBCBBCCCCCCCCCCCCCBCCCCCCCCCCCBCBCCCCBCCBCBCCCCCCCCCCCCBBBAAA9877765543322020222334555678889ABBBCCCCCCCCCCBA8644579ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBA9998887777655554443322222020000000000000335577889ABBCCCCCCCECCCCCCCCCCCCCCCCCCCCCCCCC77777777777777777776656666777777777777788888888898989899999999A9A9A9AAAAAABAABABAAABABBABABBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBBBCBCCBCBBCCCCCCCCCCCCCBCCCCCCCCCCCBCBCCCCBCCBCBCCCCCCCCCCCCBBBAAA9877765543322020222334555678889ABBBCCCCCCCCCCBA8644579ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBA9998887777655554443322222020000000000000335577889ABBCCCCCCCECCCCCCCCCCCCCCCCCCCCCCCCC;
		rom_data[507] <= 3840'h77777777777666666777777777777778888889898998998999999A9A9AAAAAAAAAAAAAAAABBBBBBBBBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBBBBBBBCCCCBCCCCCBCBCCCCCCCCCCCCBCBCBCBCCCCCCCCCCCCCCCCCBCBCCCCCCBCBBBA99887765543322202222334555778899AABBBCCCCCCCCCCCB9754578ABBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBAA9988777766555544333222220000000000000023456789AABBCCCCCCECCCCCECCECCECECCECCCCCCCCCCCC7777777777777777777666666777777777777778888889898998998999999A9A9AAAAAAAAAAAAAAAABBBBBBBBBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBBBBBBBCCCCBCCCCCBCBCCCCCCCCCCCCBCBCBCBCCCCCCCCCCCCCCCCCBCBCCCCCCBCBBBA99887765543322202222334555778899AABBBCCCCCCCCCCCB9754578ABBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBAA9988777766555544333222220000000000000023456789AABBCCCCCCECCCCCECCECCECECCECCCCCCCCCCCC;
		rom_data[508] <= 3840'h77777777777766666677777777777788888888889889999999999999A9AAAAAAAAAABABABABBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBBBBBBCCBBCBCCCCCCCCBCBBCBCCCCCCCCBCBCCCCCBCCCCCCCCCCCCCCCCCCBBBA99888765543322202223334556778899AABBCCCCCCCCCCCCCBA8544689BCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBAAA9988877766555544333322222000000000000223456788ABBCCCCCCCCCCCECCECCCCCCCCCCCCCCCCCCECCCCCC7777777777777777777766666677777777777788888888889889999999999999A9AAAAAAAAAABABABABBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBBBBBBCCBBCBCCCCCCCCBCBBCBCCCCCCCCBCBCCCCCBCCCCCCCCCCCCCCCCCCBBBA99888765543322202223334556778899AABBCCCCCCCCCCCCCBA8544689BCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBAAA9988877766555544333322222000000000000223456788ABBCCCCCCCCCCCECCECCCCCCCCCCCCCCCCCCECCCCCC;
		rom_data[509] <= 3840'h77777777777766667777778787777788888888898999899999999A9A9AAAAAAAAAAAAAABAABABABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCCCCCBCCCBCCCCCBCCCCCCCCCCBCCCCCCCCCCBCCCCCCCCCCCBCCCCCCCBBBBBAA9888765544322002223334556778899ABBBCCCCCCCCCCCCCCCB8744579ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAA99888777765554443333222200000000000000234567899ABCCCCCCECECECCCCCCCCCECCCECCCCCCCECCCCCCCECC7777777777777777777766667777778787777788888888898999899999999A9A9AAAAAAAAAAAAAABAABABABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCCCCCBCCCBCCCCCBCCCCCCCCCCBCCCCCCCCCCBCCCCCCCCCCCBCCCCCCCBBBBBAA9888765544322002223334556778899ABBBCCCCCCCCCCCCCCCB8744579ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAA99888777765554443333222200000000000000234567899ABCCCCCCECECECCCCCCCCCECCCECCCCCCCECCCCCCCECC;
		rom_data[510] <= 3840'h777777777777766677777778787777888888898889889999999999A9A9AAAAAAABAAABBABABABBBABAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBBCBCBBBBCCBCBCBCBBCCBCBCCBCCBCCCBCBCBCCBCCCBCCCCCCCCCCCBCCCCCCBBBAA9888775544322022223344556788899AABBCCCCCCCCCCCCCCCCBA854568ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAAA9988877776555544333322222202000000000003457789ABBCCCCCCCECCCCCCCECCECECCCCECCCCCCCCCCCCCECCCCCC77777777777777777777766677777778787777888888898889889999999999A9A9AAAAAAABAAABBABABABBBABAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBBCBCBBBBCCBCBCBCBBCCBCBCCBCCBCCCBCBCBCCBCCCBCCCCCCCCCCCBCCCCCCBBBAA9888775544322022223344556788899AABBCCCCCCCCCCCCCCCCBA854568ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAAA9988877776555544333322222202000000000003457789ABBCCCCCCCECCCCCCCECCECECCCCECCCCCCCCCCCCCECCCCCC;
		rom_data[511] <= 3840'h7777777777777667777777887778788888888889898998999999A99A9AAAAAAAAAAAAAABABBBBABBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCBBCBCBCBBCCCBCBCBCCCBCCBCCCCCCCCCCCBCCCCCCCCCCBCCCCCCCCCCCCCCCCCCBCBBAA998876554432220222334455677889AABBBCCCCCCCCCCCCCCCECCA8654589BCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBAAA9988877766555544333222222000000000000022355789ABBCCCECCECECCCECECCCCCCCCCCECCCCECCCECECCCCCCCCCCCC777777777777777777777667777777887778788888888889898998999999A99A9AAAAAAAAAAAAAABABBBBABBABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCBBCBCBCBBCCCBCBCBCCCBCCBCCCCCCCCCCCBCCCCCCCCCCBCCCCCCCCCCCCCCCCCCBCBBAA998876554432220222334455677889AABBBCCCCCCCCCCCCCCCECCA8654589BCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBAAA9988877766555544333222222000000000000022355789ABBCCCECCECECCCECECCCCCCCCCCECCCCECCCECECCCCCCCCCCCC;
		rom_data[512] <= 3840'h77777777777776767777788888878788888888889898989999999999A9A9AAAAAABABABABABABBBBBABBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBCBCBBBBCBCCCCBCBCBCCBCCCCBCBCBCCCBCBCCBCBCCCCCCCCCCCCCCCCCCBBBBAAA988876655433220222334555777889AABBCCCCCCCCECCCCCCCCCCCC9754578ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBAAA99888877765555444333222202002000000000023456789ABCCCCECCECCCCCECCCCECECECECECCECECCCCCCCCCCECCCECECCC7777777777777777777776767777788888878788888888889898989999999999A9A9AAAAAABABABABABABBBBBABBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBCBCBBBBCBCCCCBCBCBCCBCCCCBCBCBCCCBCBCCBCBCCCCCCCCCCCCCCCCCCBBBBAAA988876655433220222334555777889AABBCCCCCCCCECCCCCCCCCCCC9754578ABCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBAAA99888877765555444333222202002000000000023456789ABCCCCECCECCCCCECCCCECECECECECCECECCCCCCCCCCECCCECECCC;
		rom_data[513] <= 3840'h777777777777776777788887878787888888888889889899999999A9A9A9AAAAAAABAAAAAABABABABBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBBCBBBCBCBCBBCBCBCCCCCCBCBCCCCCCBCCCCCCCCCCBCBCCCCCCCCCCCCCCBBBBAA988877555433220222334555778889AABBBCCCCCCCCCCCCCCCCCCCCCA8654589ABBCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAAAA99998887777666554444333222202000000000000234567899BCCCECECCCCCCECECCCECCCCCCCCCCCCCCCCCECCECCCECCCECCCCCCC77777777777777777777776777788887878787888888888889889899999999A9A9A9AAAAAAABAAAAAABABABABBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBBCBBBCBCBCBBCBCBCCCCCCBCBCCCCCCBCCCCCCCCCCBCBCCCCCCCCCCCCCCBBBBAA988877555433220222334555778889AABBBCCCCCCCCCCCCCCCCCCCCCA8654589ABBCCCCCCCCCCCCCCCCCCCCCCCCCCBBBAAAA99998887777666554444333222202000000000000234567899BCCCECECCCCCCECECCCECCCCCCCCCCCCCCCCCECCECCCECCCECCCCCCC;
		rom_data[514] <= 3840'h7777777777777777777788888878788888888888898989989999999A9A9AAAAAAAAAAAAAAABBABBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBBCBBBBCBBBCBCBCCCBCBCCBCBCCCCCCCCBCCCCCCCBCCBCBCCBCCCCCCCCCCCCBBBAAA998877554433222223334556777899AABBCCCCCCCCCCCCCCCCCECCCCCC9754578ABBCCCCCCCCCCCCCCCCCCCCCCCBBAA99998888777777665666554433322202020000000000224457889ABBCCECCECECECECCECCECCCECECECECECECECECCECCCECCCECCCCCCCCC777777777777777777777777777788888878788888888888898989989999999A9A9AAAAAAAAAAAAAAABBABBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBBCBBBBCBBBCBCBCCCBCBCCBCBCCCCCCCCBCCCCCCCBCCBCBCCBCCCCCCCCCCCCBBBAAA998877554433222223334556777899AABBCCCCCCCCCCCCCCCCCECCCCCC9754578ABBCCCCCCCCCCCCCCCCCCCCCCCBBAA99998888777777665666554433322202020000000000224457889ABBCCECCECECECECCECCECCCECECECECECECECECCECCCECCCECCCCCCCCC;
		rom_data[515] <= 3840'h77777777777777677778888887788888888888889898989899999999A9A9A9AAAABABBBBABABBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBCBCBCBCBBCBCCBCCBCCCCCCCBCBCBCCCCBCBCBCCCCCCCCCCCCCCCCCCCCCBBBBAA998877655433222223344556778899AABBCCCCCCCCCCCECCCCCCCCECCCCA8654579ACCCCCCCCCCCCCCCCCCCCCBBAAA8888887777666665555556554323222000000000000023456789ABCCCCCCCCECCCCECCECCCECCECCCCCCCCCCCCCCCCCECCCECCECCCECECECCC7777777777777777777777677778888887788888888888889898989899999999A9A9A9AAAABABBBBABABBBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBCBCBCBCBBCBCCBCCBCCCCCCCBCBCBCCCCBCBCBCCCCCCCCCCCCCCCCCCCCCBBBBAA998877655433222223344556778899AABBCCCCCCCCCCCECCCCCCCCECCCCA8654579ACCCCCCCCCCCCCCCCCCCCCBBAAA8888887777666665555556554323222000000000000023456789ABCCCCCCCCECCCCECCECCCECCECCCCCCCCCCCCCCCCCECCCECCECCCECECECCC;
		rom_data[516] <= 3840'h777777777777777777778888888778888888888889889899999999A9A9AAAAAAAAAAAAAABABBABBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBBBCBCBCCBCBCBCCBCCCBCBCCCCCCBCBCCCCBCBCCCCCCBCCCCCCCCCCBCBBBBAA998877655433222222334556778899ABBBCCCCCCCCCCCCCCECCECCCCCCCCB9744568ACCCCCCCCCCCCCBCCCBBBAAA9887765655555555555544455543322200200000000023456789ABCCCCCECECECCECECCECCCECCCCCECECECECECCECECECCCECCCCCCECCCCCCCCC77777777777777777777777777778888888778888888888889889899999999A9A9AAAAAAAAAAAAAABABBABBBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBBBCBCBCCBCBCBCCBCCCBCBCCCCCCBCBCCCCBCBCCCCCCBCCCCCCCCCCBCBBBBAA998877655433222222334556778899ABBBCCCCCCCCCCCCCCECCECCCCCCCCB9744568ACCCCCCCCCCCCCBCCCBBBAAA9887765655555555555544455543322200200000000023456789ABCCCCCECECECCECECCECCCECCCCCECECECECECCECECECCCECCCCCCECCCCCCCCC;
		rom_data[517] <= 3840'h777777777777777777788888887788888888888898989989999999A9A9AAAAAAAAAAAABAAABBBBABBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBBBBBBCBBCBCBCBCBCCBCCCCCCBCBCBCBCCCCCCBCCCBCCCBCBCCCCCCCCCCCCBBBBBAA988877655433222223344556778899ABBBCCCCCCCCCCCCCCCCCCCCCCCCCECCA8544589BCCCCCCCCCCBA9AAAA999888766555545444444444433344433222000000000000345678AABCCCECECCCECCCECCCCECCECCECECECCCCCCCCCCECCCCCCECCCECECCCCECECCCEC77777777777777777777777777788888887788888888888898989989999999A9A9AAAAAAAAAAAABAAABBBBABBBBABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBBBBBBCBBCBCBCBCBCCBCCCCCCBCBCBCBCCCCCCBCCCBCCCBCBCCCCCCCCCCCCBBBBBAA988877655433222223344556778899ABBBCCCCCCCCCCCCCCCCCCCCCCCCCECCA8544589BCCCCCCCCCCBA9AAAA999888766555545444444444433344433222000000000000345678AABCCCECECCCECCCECCCCECCECCECECECCCCCCCCCCECCCCCCECCCECECCCCECECCCEC;
		rom_data[518] <= 3840'h77777777777777777777888887878788888888888889898899999999A9AAAAAAAAAABAAABBABABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBCBBCBBCBCBCBCCBCCCBBCCCCCCCCCCCCCBCCCCCCBCCCCCCCCCCCCCCCCCBBBBA999887765543332222334455677889AABBBCCCCCCCCCCCCECCCCCCCCCCCCCCCCB8754578ABCCCCCCCCA98778888877775555444443433333333322233222200000000000345789ABBCCCECECCCECCECECCCECCECCECCCECCCECECECECECCCECECCCECCCCECECCCCCECCC7777777777777777777777777777888887878788888888888889898899999999A9AAAAAAAAAABAAABBABABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBCBBCBBCBCBCBCCBCCCBBCCCCCCCCCCCCCBCCCCCCBCCCCCCCCCCCCCCCCCBBBBA999887765543332222334455677889AABBBCCCCCCCCCCCCECCCCCCCCCCCCCCCCB8754578ABCCCCCCCCA98778888877775555444443433333333322233222200000000000345789ABBCCCECECCCECCECECCCECCECCECCCECCCECECECECECCCECECCCECCCCECECCCCCECCC;
		rom_data[519] <= 3840'h77777777777777777778888888787888888888888898889899999999A9A99AAAAAAAAABBABBBBBBBBBBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBCBCBBCBBBBBCBCCBCBCCCCBBCCCCCBCBCCCBCBCBCCBCCCCBCCCCCCCCCCBBBAA99887765543332233334455777889AABBCCCCCCCCECCCCCCCCCCCCCCECCECCCCB98544578ABBCCCCCB8755556766656555444333232222222222220222020000000002345789BCCCCECECCCCECCCECCCCECECCCCECCECCCECCCECCCCCCCECCCCCECCCECCCCCCECECCCEC7777777777777777777777777778888888787888888888888898889899999999A9A99AAAAAAAAABBABBBBBBBBBBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBCBCBBCBBBBBCBCCBCBCCCCBBCCCCCBCBCCCBCBCBCCBCCCCBCCCCCCCCCCBBBAA99887765543332233334455777889AABBCCCCCCCCECCCCCCCCCCCCCCECCECCCCB98544578ABBCCCCCB8755556766656555444333232222222222220222020000000002345789BCCCCECECCCCECCCECCCCECECCCCECCECCCECCCECCCCCCCECCCCCECCCECCCCCCECECCCEC;
		rom_data[520] <= 3840'h77777777777777777778888887877788888888888898989998999999A99AAAAAAAAAAAAABABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBCBCBBCBBBBCCBCBCBCBCCCCBCBCCCCCBCCCCCCCCCCCBCCCCCCCCBBBCBBAA98887765544322322334556777899ABBBCCCCCCECCCCCCECCCCECCECCCCCCCCCCCB87544579BBCCCCBA85434455555555544333322222202022222000000000000002346789BCCCCECECCECECCCECCECECECCECECCECECECCCECCCECECECCCECECCCECCECECECCCCCECCC7777777777777777777777777778888887877788888888888898989998999999A99AAAAAAAAAAAAABABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBCBCBBCBBBBCCBCBCBCBCCCCBCBCCCCCBCCCCCCCCCCCBCCCCCCCCBBBCBBAA98887765544322322334556777899ABBBCCCCCCECCCCCCECCCCECCECCCCCCCCCCCB87544579BBCCCCBA85434455555555544333322222202022222000000000000002346789BCCCCECECCECECCCECCECECECCECECCECECECCCECCCECECECCCECECCCECCECECECCCCCECCC;
		rom_data[521] <= 3840'h7777777777777777778888888877878888888888888898998999999999A9AAAAAAABABAABBBABABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBBBBBCBCBCBCBCBCBBCBCCCCBCCCCBCCCCCCBCCCCCBCCCCBCCBCCCCCCCCCCCBBBBA998887765543332223334555778899AABBCCCCCCCCCCCECCCCECCCCCCCECCCCCECCCBA86545689BCCCCC875334455545444433322220000000000000000000000000245678ABCCCECECCCECCCCECECCECCCCECECCCCECCECCCECCCECCCECCECECCCECECCECCCCCCECECCCEC777777777777777777777777778888888877878888888888888898998999999999A9AAAAAAABABAABBBABABBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBBBBBCBCBCBCBCBCBBCBCCCCBCCCCBCCCCCCBCCCCCBCCCCBCCBCCCCCCCCCCCBBBBA998887765543332223334555778899AABBCCCCCCCCCCCECCCCECCCCCCCECCCCCECCCBA86545689BCCCCC875334455545444433322220000000000000000000000000245678ABCCCECECCCECCCCECECCECCCCECECCCCECCECCCECCCECCCECCECECCCECECCECCCCCCECECCCEC;
		rom_data[522] <= 3840'h77777777777777777778888888877888888888898898998999999999A99A9AAAAAAAAABAABAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBCBBBCBCBCCBCCBCBCBCBCCCCBCBCCCBCBCCCCBCCBCCCCCCCCCCCCCBBBBA99887765444322232344555778899AABBBCCCCCCCECCCCECECCCECCCECCCECCCCECCCB97544578ABBCCB8655455555444443322220000000000000000000000000245678AACCCCCCECCECCECECCCCECCCCECCECCECECCECCECCECECCECCECCCCCECCCCECCECECECCCCCECCC7777777777777777777777777778888888877888888888898898998999999999A99A9AAAAAAAAABAABAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBCBBBCBCBCCBCCBCBCBCBCCCCBCBCCCBCBCCCCBCCBCCCCCCCCCCCCCBBBBA99887765444322232344555778899AABBBCCCCCCCECCCCECECCCECCCECCCECCCCECCCB97544578ABBCCB8655455555444443322220000000000000000000000000245678AACCCCCCECCECCECECCCCECCCCECCECCECECCECCECCECECCECCECCCCCECCCCECCECECECCCCCECCC;
		rom_data[523] <= 3840'h7777777777777777788888888888788888888888888889989899999999A9AAAAAAAAAAAABABBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBBBCBCBCBBBBCBBBCBCBCBCBCBCBBCBCCCCCCBCCCCCCBCCCCBCBCCCCCCCCCCCCCCCBCBBBAA99887765543322232334455778899AAABCCCCCECCCCCECCCCCCCCCCECCCECCCECCCCECBA87544578ABBCA87555555544443332220000000000000000000000000235678AACCCCECECCCECCECCECECECCECECCECCECECCECCECECCCCCECCECCECECCCECECCCCCCCCCECECCCEC767677777777777777777777788888888888788888888888888889989899999999A9AAAAAAAAAAAABABBBABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBBBCBCBCBBBBCBBBCBCBCBCBCBCBBCBCCCCCCBCCCCCCBCCCCBCBCCCCCCCCCCCCCCCBCBBBAA99887765543322232334455778899AAABCCCCCECCCCCECCCCCCCCCCECCCECCCECCCCECBA87544578ABBCA87555555544443332220000000000000000000000000235678AACCCCECECCCECCECCECECECCECECCECCECECCECCECECCCCCECCECCECECCCECECCCCCCCCCECECCCEC;
		rom_data[524] <= 3840'h7777777777777777778888888887778888888888888889898989999999A9AAAAAAAAAAAAAAABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBCBBBBCBBCBBCBCBCBCBCBBCCCCBCCCBCCCBCBCCCCCCCCCCCCCCCCCCCCCCBCBCBBBAA99887765543333222334555678899AABBCCCCCCCCCCCCCCECCECECECCCECCECCCCCCCCCCBA85445689ABA9876666555543332220000000000000000000000000024578ABCCCCECCCCCECCECCCECCCCCECCECECECECECCECECECCCECECCECCECCCCECECCCCCECECECECCCCECCC667676777777777777777777778888888887778888888888888889898989999999A9AAAAAAAAAAAAAAABBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBCBBBBCBBCBBCBCBCBCBCBBCCCCBCCCBCCCBCBCCCCCCCCCCCCCCCCCCCCCCBCBCBBBAA99887765543333222334555678899AABBCCCCCCCCCCCCCCECCECECECCCECCECCCCCCCCCCBA85445689ABA9876666555543332220000000000000000000000000024578ABCCCCECCCCCECCECCCECCCCCECCECECECECECCECECECCCECECCECCECCCCECECCCCCECECECECCCCECCC;
		rom_data[525] <= 3840'h777777777777777778888888877878888888888888889899989999999999A9AAAAAAAAAAABABBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBCBBCBBBBBBCBCBCBCBCBCCBBCBCCBCCCBCCBCCCBCCCCBCCBCCCCCCCCCBCBBBBBBAA99887765543322223334555778899AABCCCCCCCCECCECCCCCCCCCCCCCECCCECCECECECCCCCA97534578899887666554443322200000000000000000000000000035789BCCCCECCCECECCCECCECECECECCCECCCECCECCECECCECECECCCECCCECCECECCCCECECCCCCECCCEECECEC66676767777777777777777778888888877878888888888888889899989999999999A9AAAAAAAAAAABABBABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBCBBCBBBBBBCBCBCBCBCBCCBBCBCCBCCCBCCBCCCBCCCCBCCBCCCCCCCCCBCBBBBBBAA99887765543322223334555778899AABCCCCCCCCECCECCCCCCCCCCCCCECCCECCECECECCCCCA97534578899887666554443322200000000000000000000000000035789BCCCCECCCECECCCECCECECECECCCECCCECCECCECECCECECECCCECCCECCECECCCCECECCCCCECCCEECECEC;
		rom_data[526] <= 3840'h77777777777777777788888888777878888888888888888899899999999A9AAAAAAAAAAABABABBBABABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBCBBCBCBBBBBCBCBBBCBCBCBCBCBCCCCBCCCBCCBCCCCCCCBCCCCCCCCCCCCCBCBCBBBBAA999887765543322222334555778899ABBBCCCCCCCCCECCCCECECECCECECCCECCCCCCCCCCECCCCA86434567887666655543322200000000000000000000000000003589BCCCCECCCECCCCCECCECCECCCECCECCECECCECECCECCECCECCECECCECCCECCCECECCCCCECECCCECCCCCCCC7666667777777777777777777788888888777878888888888888888899899999999A9AAAAAAAAAAABABABBBABABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBCBBCBCBBBBBCBCBBBCBCBCBCBCBCCCCBCCCBCCBCCCCCCCBCCCCCCCCCCCCCBCBCBBBBAA999887765543322222334555778899ABBBCCCCCCCCCECCCCECECECCECECCCECCCCCCCCCCECCCCA86434567887666655543322200000000000000000000000000003589BCCCCECCCECCCCCECCECCECCCECCECCECECCECECCECCECCECCECECCECCCECCCECECCCCCECECCCECCCCCCCC;
		rom_data[527] <= 3840'h677777777777777778888888887778888888888888888998989999999A99AA9AAAAAAAAAABABBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBCBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBCBBCBBBBCBCBCBCBCBCCCBCBCCCCCCCCCCCCBCCCCBCCCCCCCCBCBCBBBBBAAA999887765544322222334455778899AABBCCCCCECCCCCCECECCCCCCECCCCECCCCECECECCCCCECCB9754345777655555543322200000000000000000000000000004589BCCCCCCCECCCECECCCECCECCECCECECECCECECECECECECECCECECCECECECCECCCCCCECECCCECECCECECECEC66667666677777777777777778888888887778888888888888888998989999999A99AA9AAAAAAAAAABABBBBBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBBBBCBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBCBBCBBBBCBCBCBCBCBCCCBCBCCCCCCCCCCCCBCCCCBCCCCCCCCBCBCBBBBBAAA999887765544322222334455778899AABBCCCCCECCCCCCECECCCCCCECCCCECCCCECECECCCCCECCB9754345777655555543322200000000000000000000000000004589BCCCCCCCECCCECECCCECCECCECCECECECCECECECECECECECCECECCECECECCECCCCCCECECCCECECCECECECEC;
		rom_data[528] <= 3840'h67777777777777777888888888888788888888888888889999899999999999A9AAAAAAAAABABBBABABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBCBCBBCBBBBCBBBBBBBCBBCBCBCBCBCBCBCBCCBCBCCBCCCCCCBCBCCCBCBCBCBCBBBBBBAAAA999887765543332222334455778899AABBCCCCCCCCECCECCCCCCECECCCCECCCCECCCCCCCECECCCCBA8543455655555554332200000000000000000000000000000358ACCCCCECECCCECECCCECCECCCECECCECCECECCECECCECCECCECCECCECCCCECECECECECCCCCECCCCECCCCCCCCC6666676667777777777777777888888888888788888888888888889999899999999999A9AAAAAAAAABABBBABABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBCBCBBCBBBBCBBBBBBBCBBCBCBCBCBCBCBCBCCBCBCCBCCCCCCBCBCCCBCBCBCBCBBBBBBAAAA999887765543332222334455778899AABBCCCCCCCCECCECCCCCCECECCCCECCCCECCCCCCCECECCCCBA8543455655555554332200000000000000000000000000000358ACCCCCECECCCECECCCECCECCCECECCECCECECCECECCECCECCECCECCECCCCECECECECECCCCCECCCCECCCCCCCCC;
		rom_data[529] <= 3840'h66676777777777777888888888888888888888888988898899998999999A9AA9AAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBBBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBCBBBCBCBBCBBBBCBCBCBCBCCCCCBCCCCCBCCCCCCCCCCCBCCBCBCBBBBBBBAAAA9988887765544332222333455778889ABBBCCCCECECCCCECCECECECCCCECECCECECCCECECCCCCCECECB9754555655555443320000000022222000000000000000002579BCCECECCCCECCCCCECCCECCECECECECCECCECECCECECCECCECECCECECECECCECCCCECCECECCCECECCECECECEC6666666666676777777777777888888888888888888888888988898899998999999A9AA9AAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBBBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBCBBBCBCBBCBBBBCBCBCBCBCCCCCBCCCCCBCCCCCCCCCCCBCCBCBCBBBBBBBAAAA9988887765544332222333455778889ABBBCCCCECECCCCECCECECECCCCECECCECECCCECECCCCCCECECB9754555655555443320000000022222000000000000000002579BCCECECCCCECCCCCECCCECCECECECECCECCECECCECECCECCECECCECECECECCECCCCECCECECCCECECCECECECEC;
		rom_data[530] <= 3840'h66667677777777777888888888888888888988889889889989899999999999A9AAAAAAAABAAABABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBBBBBBBBBBBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBCBBBBBBBBBBBBBCBBCBCBBCBCBBBCCBCCCCCCCBCCBCCCCCCCCCCCBBBBBBBAAA99888877665543322222234455778899ABBBCCCCCCCCCCECCCCCCCCCCCECCCCECCCCCECCCCECECECCCCCCA87555666555543322000002344333220000000000000000359BCECCCCCCECCECECECCECCCECCECCCECECCECCECECCCECECECCECECECCCCECECECECCECECCECECCCECCCCECCEC6666666666667677777777777888888888888888888988889889889989899999999999A9AAAAAAAABAAABABBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBBBBBBBBBBBBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBCBBBBBBBBBBBBBCBBCBCBBCBCBBBCCBCCCCCCCBCCBCCCCCCCCCCCBBBBBBBAAA99888877665543322222234455778899ABBBCCCCCCCCCCECCCCCCCCCCCECCCCECCCCCECCCCECECECCCCCCA87555666555543322000002344333220000000000000000359BCECCCCCCECCECECECCECCCECCECCCECECCECCECECCCECECECCECECECCCCECECECECCECECCECECCCECCCCECCEC;
		rom_data[531] <= 3840'h666667777777777777888888888888888888888989889989998999999999A9A9AAAAAAAAAAABABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBBBBBBCBBCBCBBCBCBCCCBCCCBCBCCCCCCCCCCCBCBCBBBBBBAAAAA9988888776655433322222344456778899ABCCCCCECECECECCECCCECECECCCECCCCECCECCECCCCCCCCECECCB8866666555443322000024565543322200000000002000247ABCCCECECECCECCCCCCECCECCCECCECCECECECECCECECECCECCECECCCECECCECCECECECCECCCCCCECCCECECCECC66566666666667777777777777888888888888888888888989889989998999999999A9A9AAAAAAAAAAABABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBCBCBBBBBBCBBCBCBBCBCBCCCBCCCBCBCCCCCCCCCCCBCBCBBBBBBAAAAA9988888776655433322222344456778899ABCCCCCECECECECCECCCECECECCCECCCCECCECCECCCCCCCCECECCB8866666555443322000024565543322200000000002000247ABCCCECECECCECCCCCCECCECCCECCECCECECECECCECECECCECCECECCCECECCECCECECECCECCCCCCECCCECECCECC;
		rom_data[532] <= 3840'h6666667777667677777888888888888888888989989989989999999999999A9A99AAAAAAABAABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBCBBCBBCBCBBBBBBBBBBBCBCBBBBBBCBCBCBCBCBBCBBCCCCCBCBCBCCBCBCBBBCBBBBAA9A9998888776655444322222233455677889AABBCCCECCCCCCCCCCCCECCCCCCCECCECECCECCCCCCCECECECCCCCCA8877775555433220002345777543220000002022220202358BCCECCCCCCCCCECECECCECCECECECECECCECCECCECCECCECCECECECECCECECCECCECCECECECECECCECECCCECCEC566556666666667777667677777888888888888888888989989989989999999999999A9A99AAAAAAABAABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBCBBCBBCBCBBBBBBBBBBBCBCBBBBBBCBCBCBCBCBBCBBCCCCCBCBCBCCBCBCBBBCBBBBAA9A9998888776655444322222233455677889AABBCCCECCCCCCCCCCCCECCCCCCCECCECECCECCCCCCCECECECCCCCCA8877775555433220002345777543220000002022220202358BCCECCCCCCCCCECECECCECCECECECECECCECCECCECCECCECCECECECECCECECCECCECCECECECECECCECECCCECCEC;
		rom_data[533] <= 3840'h56566667667667777778788888878888888889898989899999999999999A9A99AAAAAAAAAAABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBCBCBCBCBCBBBBBCBCBCBCBBBCBCBCCCCCBCBCBCCCCCCBBCBBBBBBBAAA9A99988888776655543332202233455577889AABBCCCCCCECECECECECECCECECECCCECCCCECCECECECCCCCCCECCCA98767776554432200023557887532000222222220202224579CCCCCECECECECCCCCCCECCECCECCECCECECCECCECECCECCECCECCECECECECECECECCECCECCCCCCCECCCCECCCECC6656665656566667667667777778788888878888888889898989899999999999999A9A99AAAAAAAAAAABBBBBBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBCBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBBBBCBCBCBCBCBBBBBCBCBCBCBBBCBCBCCCCCBCBCBCCCCCCBBCBBBBBBBAAA9A99988888776655543332202233455577889AABBCCCCCCECECECECECECCECECECCCECCCCECCECECECCCCCCCECCCA98767776554432200023557887532000222222220202224579CCCCCECECECECCCCCCCECCECCECCECCECECCECCECECCECCECCECCECECECECECECECCECCECCCCCCCECCCCECCCECC;
		rom_data[534] <= 3840'h656666667767667777788888888787888888889889899999999999999999999A99AAAAAAAABABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCBBBCBBBBBCBBBBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCCBCBCBBBBBCBCCCCCCCCCBCBCBCBBBBABAA99998888877665554433322222334556778899ABBBCCCCCCCCCCCCCCCCCECCCCCCCECCCCECCCCCCCCCCECECECCCB987666676555432200022457787542000002222222220224579BCECECCCCCCCCCECECECCECCECCECCECCECCECECECECECECECECECECECECCCCECCCECECECCECECECCCCECCCECCEC56565565656666667767667777788888888787888888889889899999999999999999999A99AAAAAAAABABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCBBBCBBBBBCBBBBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBCBCCBCBCBBBBBCBCCCCCCCCCBCBCBCBBBBABAA99998888877665554433322222334556778899ABBBCCCCCCCCCCCCCCCCCECCCCCCCECCCCECCCCCCCCCCECECECCCB987666676555432200022457787542000002222222220224579BCECECCCCCCCCCECECECCECCECCECCECCECCECECECECECECECECECECECECCCCECCCECECECCECECECCCCECCCECCEC;
		rom_data[535] <= 3840'h5565666676676777777878788787878888888888989898999999999999AA9A9A9AAAAAAAABABAABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCCBBBBCBBBBBBBBCCBCBBCBCBBCBCCBCCCBCBCBCBCCBBBBBBBAAA999888888777655544433322222334455778899ABBBCCCCECECECECECECECCCECECECCCECECCECECECECECCCCCCCB87555555555543320000234566654220000222322220022368ABCCCCCCECECECECCCECCECCECCECECECECCECECCECCCECECECECECCECCECECECCECECCCECCECECECCECECCECCCECC556555555565666676676777777878788787878888888888989898999999999999AA9A9A9AAAAAAAABABAABBBABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBCBBCBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCCBBBBCBBBBBBBBCCBCBBCBCBBCBCCBCCCBCBCBCBCCBBBBBBBAAA999888888777655544433322222334455778899ABBBCCCCECECECECECECECCCECECECCCECECCECECECECECCCCCCCB87555555555543320000234566654220000222322220022368ABCCCCCCECECECECCCECCECCECCECECECECCECECCECCCECECECECECCECCECECECCECECCCECCECECECCECECCECCCECC;
		rom_data[536] <= 3840'h5556566676666677777777787877788888888888888889899999999999A9A9A9AAAAAAAAABAABBAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBBBBCBCBCBBCBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBCBBCCBBCBCCBCBCCCCBCCCBCCCBCBCBCBBBBBBBBAA999888877776655444333222022333455678899ABBCCCCECCCCCCCCCCCCCCCECCCCCCECECCCECCCCCCCCCCECECCCA854445554444442200000023444432200000022222222002589BCCCCCECCCCCCCCCECCECCECCECCECCECCECECCECECECCECECCECCECECECCECECECCECECCECECECCECECCECECECCEC555555555556566676666677777777787877788888888888888889899999999999A9A9A9AAAAAAAAABAABBAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBBCBBBBCBCBCBBCBBBBCBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBBCBBCCBBCBCCBCBCCCCBCCCBCCCBCBCBCBBBBBBBBAA999888877776655444333222022333455678899ABBCCCCECCCCCCCCCCCCCCCECCCCCCECECCCECCCCCCCCCCECECCCA854445554444442200000023444432200000022222222002589BCCCCCECCCCCCCCCECCECCECCECCECCECCECECCECECECCECECCECCECECECCECECECCECECCECECECCECECCECECECCEC;
		rom_data[537] <= 3840'h55656666667676777777878777777788888888888888988999999999999A9A9A9AAAAAAAAAABAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBCCBCBCBBCBCCBBCCBCBBCBCBCBCCBCBCCBBCBCBBCBBAAAAAA9998888777665554443332222022233455678899AABCCCCCCCECECECECECECECCCECECECCCCECCCECECECECCCECBA8753235555433323200000002333323220200002222220222368BCCECCECCECECECECCCECCECCECECCECCECECCECCECCECECCECECECECECECECCECCECCECECCECCCECECCECCCCECCECC5555555555656666667676777777878777777788888888888888988999999999999A9A9A9AAAAAAAAAABAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBCCBCBCBBCBCCBBCCBCBBCBCBCBCCBCBCCBBCBCBBCBBAAAAAA9998888777665554443332222022233455678899AABCCCCCCCECECECECECECECCCECECECCCCECCCECECECECCCECBA8753235555433323200000002333323220200002222220222368BCCECCECCECECECECCCECCECCECECCECCECECCECCECCECECCECECECECECECECCECCECCECECCECCCECECCECCCCECCECC;
		rom_data[538] <= 3840'h656566666667676777777777777777788888888888888888989899999A99A9A9AAAAAAAAAAAABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCCBBCBCBBBCCBCBCCBCBCBCCCBCBCCCBCBBCBBBABAAAAA9998887777655554433322220222233455678889ABBBCCCCCCCCCCCCCCCCCCCCCECCCCCCCCECCCECCCCCCCCCECCB975332235655422220200000002222222220000020222220202379BCCCECCECCCCCCCCCECCECCECCCCECCECECCECCECCECECCECECECCECCECCECECCECECECCCECCCECCCCECCCECECECCEC55555555656566666667676777777777777777788888888888888888989899999A99A9A9AAAAAAAAAAAABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBCBCCBBCBCBBBCCBCBCCBCBCBCCCBCBCCCBCBBCBBBABAAAAA9998887777655554433322220222233455678889ABBBCCCCCCCCCCCCCCCCCCCCCECCCCCCCCECCCECCCCCCCCCECCB975332235655422220200000002222222220000020222220202379BCCCECCECCCCCCCCCECCECCECCCCECCECECCECCECCECECCECECECCECCECCECECCECECECCCECCCECCCCECCCECECECCEC;
		rom_data[539] <= 3840'h66566666667667677777777777777778888888888888888889898999999A9A9A9AAAAAAAAAAAABABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCCCCBCBCBCBCBCBCCBCCCCBCBCBBBBBBABAAA999998887776555554433222220202233455677899AABBCCCCCCECECECECECECECECCECECECECCCECCCECECECECCCB9743223345554322000200000000222222000202022222202022579CCCCCCECCECECECECCCECCCCCECCECECCCCECCECCECCCECCECCCECCECCCECCCECECCECECECCECECECECCECCCCCCCECC5555555566566666667667677777777777777778888888888888888889898999999A9A9A9AAAAAAAAAAAABABBABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCBBBCBBCCCCBCBCBCBCBCBCCBCCCCBCBCBBBBBBABAAA999998887776555554433222220202233455677899AABBCCCCCCECECECECECECECECCECECECECCCECCCECECECECCCB9743223345554322000200000000222222000202022222202022579CCCCCCECCECECECECCCECCCCCECCECECCCCECCECCECCCECCECCCECCECCCECCCECECCECECECCECECECECCECCCCCCCECC;
	end
	
	// =======================================================
	// Data
	// =======================================================
	reg		[10 : 0]		rom_y;
	reg		[3839 : 0]		tmp_data;
	
	wire	[lut_bw*2-1 : 0]		data_t0;
	wire	[lut_bw*2-1 : 0]		data_t1;
	wire	[lut_bw*2-1 : 0]		data_t2;
	wire	[lut_bw*2-1 : 0]		data_t3;
	
	assign data_t0 = gray_lut[tmp_data[3839 : 3836]] << {gray_cmp, 1'b0};
	assign data_t1 = gray_lut[tmp_data[3835 : 3832]] << {gray_cmp, 1'b0};
	assign data_t2 = gray_lut[tmp_data[3831 : 3828]] << {gray_cmp, 1'b0};
	assign data_t3 = gray_lut[tmp_data[3827 : 3824]] << {gray_cmp, 1'b0};
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			
			epp_data_r <= 8'b1010_1010;
			rom_y <= 11'd0;
		end else if(
			(cnt_b >= (fsl + fbl - 1)) &&
			(cnt_b < (fsl + fbl + fdl - 1))
		)begin
			if(
				(cnt_a >= (lsl + lbl - 1)) && 
				(cnt_a < (lsl + lbl + ldl - 1))
			)begin
				
				if(disp_all_w)begin
					epp_data_r <= 8'b1010_1010;
				end else if(disp_all_b)begin
					epp_data_r <= 8'b0101_0101;
				end else begin
					// epp_data_r[15:14] <= tmp_data[0] ? 2'b10 : 2'b01;
					// epp_data_r[13:12] <= tmp_data[1] ? 2'b10 : 2'b01;
					// epp_data_r[11:10] <= tmp_data[2] ? 2'b10 : 2'b01;
					// epp_data_r[ 9: 8] <= tmp_data[3] ? 2'b10 : 2'b01;
					epp_data_r[ 7: 6] <= data_t0[lut_bw*2-1 : lut_bw*2-2];
					epp_data_r[ 5: 4] <= data_t1[lut_bw*2-1 : lut_bw*2-2];
					epp_data_r[ 3: 2] <= data_t2[lut_bw*2-1 : lut_bw*2-2];
					epp_data_r[ 1: 0] <= data_t3[lut_bw*2-1 : lut_bw*2-2];
				end
				
				tmp_data <= {tmp_data[0+:(3840-4*4)], 16'd0};
			end
			
			if((cnt_a == (lsl + lbl - 1 - 1)))begin
				tmp_data <= rom_data[rom_y];
			end
			
			if(cnt_a == (lsl + lbl + ldl - 1))begin
				if(rom_y >= (540-1) )begin
					rom_y <= 11'd0;
				end else begin
					rom_y <= rom_y + 1'b1;
				end
			end
		end
	end
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			gdck_r <= 1'b0;
		end else begin
			if(
				(cnt_a >= (lsl + gdck_sta - 1)) && 
				(cnt_a < (lsl + gdck_sta + gdck_hi - 1))
			)begin
				gdck_r <= 1'b1;
			end else begin
				gdck_r <= 1'b0;
			end
		end
	end
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			gdsp_r <= 1'b0;
		end else if(cnt_a >= (ltot - 1))begin
			if( cnt_b <= (fsl - 1) )begin
				gdsp_r <= 1'b0;
			end else begin
				gdsp_r <= 1'b1;
			end
		end
	end
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			sdoe_r <= 1'b0;
		end else if(cnt_a >= (ltot - 1))begin
			if(
				(cnt_b >= (fsl + fbl - 1)) &&
				(cnt_b < (fsl + fbl + fdl - 1))
			)begin
				sdoe_r <= 1'b1;
			end else begin
				sdoe_r <= 1'b0;
			end
		end
	end
	
	always@(posedge glb_clk)begin
		
		if(!glb_nrst)begin
			gdoe_r <= 1'b0;
		end else if(cnt_a >= (ltot - 1))begin
			if(
				(cnt_b >= (fsl - 1)) &&
				(cnt_b < (fsl + fbl + fdl - 1))
			)begin
				gdoe_r <= 1'b1;
			end else begin
				gdoe_r <= 1'b0;
			end
		end
	end
	
endmodule
